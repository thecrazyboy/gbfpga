��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�ϗ7�#���H�����u�g[iˬ���t|�3���ҥ�ys�B�@Yq�"F}�\"QY����#�ڇ7�\ӷ��繟��1W�k���q�u ���{�m)RM�S|@�����ͣz��yʿG��O�Yg>�s$h_!��-~���=wx�=�M�����/�mb�K#�� ��1��W�i�{,?�EM�N�0�K
䧣�:39ok^�(��-���V�f���Sk�	����}ؖŸ�*����~������6l@ޱ����t����_.��±7�Eۨ[�ܐb\T�8�����"��!'���^C�he�K�Zw��J�;��E���a�BnB��lje8�i�U��^w�K�@ܚ��^<'�������������a}��a��W��S��!�P�:�ޓ��|=ǎO�k�σf&�_ K(yǦ�+F{v5�X�x!}e�y�D��"љn3]��6:�Ѳ=&:_��h�,�klf�es�4�=|��-�#3��r�E8m>�e7�{�~w���O3��{	 X�n���7��[��{d�mҫFG�6�ݝZ���4́���GF��yw�D��Օ��挹O����[�K6���L���ڹ�\Z'�
���lS}d}��w7�� ^$�j_��묡X<P�`��&X���xRq�y��G���R��B�}[�b50t��j�k\��Ju�a�V�ؒ���w�\%RF�Z�購�:*EO�GT+���,��B�/�9K�5J���t	���y"q��yǕR�<�]���>{�t�f�'z�(*��l�����'J|N�]�F����Yz�ȅy��/��)�B��
�vu`o9M5|�Z�e������gM"���C�W��f,�o�`��<��Xk�:�s#�T��/q�PC���k�!}5������j��b%׊a1-�b��\%猢��S������Ew�Z���UYwds�i��;�IT'q��z9}j��!/m�n��4�Z������ء�\��0d��>�fZ{�>�Q���}o�x�/=̪Y�I�s<T�y-���G���_�җ���2���5�g�$K�+�'y��wj�%��� ����s�ٸe�p{��V�$C؄��G��Q}����P�fr#ZY_.&;�i�[!CY�V�B�s͓8�ճx��L�[s��́;��U,�������_�sԫ��խ�[)Hc�F��
�ɂ�I;1l�T;�n���:5z�P_=#�M$�.��O���q�'��1 BO�>�%���p�3_���T�����s����~A���A�}��[�x��SwT A½�Nn�&��!��I) ���`� ���QH����;�b���f��zJ���(�����s�C�'l��HC�j���	�ajG������D�s�C���<�L&<p��໧���l��x8u����^p�/}8#C���v����<����ʪ���)�#��4���LL�g۹�N����$]��$T�3<�Q�Wؾ�	���~���Nmؼ*q^��$���r�h� ѣ�|x�OM��o!�j	?�Zm�.x�����o�
��xKH$�Ni4�CjˋzV>��gD~�T����Ec��$(�̽����I ��r:!���іm�*�m�d�YIj�y54~HD�jZ5�� .�k���^��x����k*�0��A�C[AiZS���y4�!l�T(G�Q(h;g��?V�eA�H�2���s�?�f�S�Ln|��<���Q9��N��L��']��5⊭��'���w��Q����o���)�A3�(m�k89����%(k������)�3Kg<�{X[�j�����˨V�XnXI>�ֻ;�,s-�+���x�5qRL�s�=�Ɵ�|H��e\��[�g����l���p�kq2��X�V*�	��u{�Q�5M�8>{�꣣��bJe#x0Ul.H;܄�	��_N`J(v�{�u�%*�J!apyÜEr��'k-���W������qJy��I���$��	��ɢ�����f��侳������#B���a����.:"01��Kp~�~�,t��M�0Yo�����)�F`�/]!��0�13������y�y!�$tNYp�?Y� #M&�m�b��B��.��� ��"p���Գ_���/�:�SD�w���^�K��:�����rѨ�l�!ȳ����XP<V�5���F�!O ЗkΆ�������@U�(��������5�<1�qY�bB�8(���,	G���ٷ'��b��
�X�Z
{L&�6"'�j�Z&9���3`��OЗ��,��?�U��L��W��d��0}CV� le�o4q�tSJ|c�i�"D����⏜���V!���c]����S�|2����z���U�+������kO�n0�o����+#�"v��]��YɁFK�&rѹn��S������m7��ĘB�{�\��`d����Ʋ6�^�ړ*��ް�.w��~B �Yi��;R�I����Ǽ=5zy�:�(�o+��5]P��\1WZ2�&G�I�\KHB2�V�Ğ�ozrz�5G�k�(Z��R�:P0s5#��q��/U��b�t�ۜ`SC�fE~��2�p*���ʘ#�`T'��x��7���9�g}}��W�B�f��"�.��~ކ�FI![Ur>�г�t�k���-So�g?dX@nA�G����T���:�+I�}�{��� �̜Mz��ܹ�I8�V��*9o�����������5Ӎ�E�M�$�S~vsČ]{�B�̊08kj:1�)�*_�s��eΥ�)d�
�L�fpw9�-m6��mG:ݥg�2�M�(�Bn?� "R׉����.#{��pX��$�'o�n3�i�E����'���)P�&�����_�Y���
J�����U4����n
c��V��0R���u3�s�/'������?��i��"�	���!��Ҿ������ i>�tydZ�%ϳ��}��K	�"(�ߠ}ax+����?({얍gU�����%��q)�[yM�V��)F �ZCK8J�B�k��Ѵ�K�[_nP�}��������]ؙɄЛ��зJ�}�$du-[P��ޯ�Φ3��H~�a�t��P�]�T��llZ&�!O�#&ݺ�YӔE�]X�6-�1�b��u\#0�8֍9��@S��o�����i�N��X��ɸ<��}^t�Lp�H��چJ�a��?�J��@-q E�sf��;�r;Ze�q��������j�	͜���[���҂��^B��{+��޹'�:�)?��I���ټ�}��Tԋ�4:%�|8NGʊ��L��o�U�?���u���q*��3� ������t��Th�*Z��n���C/���U����(P��kB>�>��[x���H5��Z-�q�"^�+��<���R	����	z��(9%ܸ�b\��_����Ӣ$�_���#扱N�\B�T4f����r~%��Q00ҟ,��z���ܕ���ռ�+�/U�`2 a�SzDemS	U;��C2�vQL�ȿ]ծ��$89ҧ�]�������Vc�JUi�̴����1�ʞ��G��,�3i%I'�$l��i�w�%�3�\NyH�%L�_�G��Q���.��D�B����1�A�RU�~��|��W����>ŏ6�/>��+Tg�|�f����Y��U�ƥ�� ���	��wm���
ӝ"��/����>��!B����eP�{M[+B�UTy���b�!�W�Ѧ��ԝ1�VK�������R���w��'9�s����-?]����$�{b��id�R�6/�k��7
%�JYmãz#���d�=,3���`��1��	�+'��a?�DÀ�?�6�{�QC��+�`�� ��
��Z���X��mx�ZR�;���d;R�{n���J�S�N+������Oܩqy����w�3�e�4�BxU)�(.�RE�$#~b��'�_N�������}ty���^s�83��-�R>ڂ|�U�8�VWM�y�m�a���C�ޯ����)�P���;�s~p)f�~1+�.g��(�s�u`� ���ԂǸe�@��+=��i���IaމI�ը\Ƃ/�_���Ԡ;���7�O�0I.����N���S��5/�BoO���΂`97B�L�%������V�~R`Ȱ�:��Qg ���m�A�����j�ӊ����ӳ��ފ᪉�=�c�λ��RK�����g�67%��y��	̻~���{2��,�?�d("�ERi�V>��R�xr�@)А\�i�_��ZR��AlWw,�z��G<o���;#Z�Q�@�A*!�]��	tt1�d����¦N+�P��hgJ��m��n%Sw�^
 ;�ȥ�&ɟ�u�$�VJ���T��\� �Px�6�+F0V���!��e`�ާ��/�����%~�g�����Ͼa�o�;�7؊}����RV'��U*����̐�wܵ��7+
�;ϚЊ��0r)�:C�/���SݼOFB�^.f�IM��pL����ZF:���"��bJ�.�%����*�J^c �]�l�Z��f�i���(�|8��0�l�c�[���ܶ ���E�Z��@Ӛ����;�`�k�yo�NȄwOƻ7�̈́��"�u�
�������ׁ�����/��"�Iߞ"zuOv;_~��d��:ȴ�y9�c]ˡc@�m�ȀR���:YR}�����1��IH����/=�`q	!p�wXU��D85̀PYL�ضݷG��X0U��-��� �h�T>:b(�=o���GZ��Ҭ��dK��4S;E�Uz����Ju��O%��`��~�X��*����d4�5�G�9Μ ����LsWs��( N{�R�mw^5�>���C�����S�U�1���OS��ߏ��'\q*�h<��=�kSF"�+�����5�ج������j?��ֆ^�f${�P��C��R���_�o��B=�тCq��Y��{���� �u=z=�:9I �����mX�o9P)�5S"�l^ݻ���TόRl��Z��i��Gr/�D�ˆ��s!���uC���k�H�ç�0Vc�<Qx�y�Y��D�k�9
'��sHV@Jp������B'7�p͌;b���=)�%}n	�E���W�;�r:�\�rJP}w���Ga��Cכ������%4�	>��!y�������^I�J�2�g�é^�ʃ}L�1=�w�p�|b/���4�+>�u?�]�W��(-0Dnq�B�%Lk쪵7�n=Q�B#uF��D�������a���)��)��_�5�����<M�&��9b┎���vOl�i,��LM&�}JL4Ѻ3?�5/Y����8�>|+dU�� w�H�T�p��+i�ҧ�//��T�C�4��_�u�l�k�34�
z/�_Av�db@e������t��<�=�`�3zFq(6��7>�> \݁��,^~-�7�Ν�q�{n���L}���E-9�-!����Ԉ�:6�g��7�(4�R{��!eB�����W���';��*h��Q����w�c���\t�.E��^�&*���Qٮ=��n�j���	�Dp_��Aoƾ�t<��W����B�X�z.2��뿗�AP�!c�@��[ָ9�E��ܐ�?������M�!)�2���t>�KaO<G�X���w�hO��oP��>c҈%�[���#lQ쭱:� �õ�Z�(�B5���7�SQ�V�6Bh�ʗ_Nt�V9ܫ�t��	mo�I6,Z������Ӿ=����QsW���(��ߚm�TgΎ�Ւ��!؃z��W���//Pw�;��V��!@��|����n=��2��=�gBNo\���E�����x���r�kw��s��ޫ��0vf�^����܎�G2_�ҾuH���i��V�X�؜o���;0�� �/������>$n��JA�����#�zWSt�0(}��d����\ld�5�c��wj)�
�Q��qtt]�;�DG�5)4��ձn��׫�A�ׇ�o��Xb&q�I�W�uF�U+P���:�W?O��'�">`.�~P��2���[q�"�>	�y��"�����V>��#����t�m�,�l
��R���H�I�;T�(�q�E�-���@cc�8�I��7p�u�/ܾ�)��͈!�KA�$�+� ><�}��ؿ��O�r\��/������o��b��$uci�b�e-
~zӒb�?_�K��|Hi���L�Ԓ�Ƶ�1n��nT,����hqp���2���ezPVIb��W:���e�U��C ���];Sa>����������͟p5���a�B�����Lo��yv�p(��=��|��8��,�A��8�8���[Z�i����n�ngp���\��=��K'�!���[ eT�&	ʶ,����q���pz�Ψ����hO���p��q��n%8}O�S+��5=K9
�H��I�Ŀ�t���+��F�|C�Դv�``�����N�9��Z$O܅X��&��C�/W�M@"1�LN�6��{W�i�;�o�20�7�o1�>1C7n�k~�]2�^|�ճ����\�������'iT��V�i�zZRI���0z�-���qU���2~*�ğP����15�yW�����G��Q���h� D>�l�g��&��u,ρ�����e9�U�&��t?��c=����Y�p|�)Fd7����~/��'~��
p�X�C�'p4uL��m����_)-^�m2Q(RU�O(�T��}�"��07��"��k·� /�����U�,�ᣁ�Ъ��N�غB�sY"ƆaW�6�O5aQ�<�%@��@R������h��� ��qsn���u2_!��cBܞ~��ɯ%�'�����Yzx��3c�ʌmt�V �$O7 ��D@ꭤ鶕��u���z��h�[�"Y��:����!Cp�g�
R���T�H���k�V�M�C�ٝ�M��q8�_#�D,��,ڐ��ȈV4r��A����1��gџ�:ޠk���e�(���2;�z�ۙ�0�	�M}ֱA-X`���zM�yvHQ�s�o�B���m]x�î	�1X��)���#��Yd���o���K�:\}dN>�!��W{y�,)�ʧ{w�%Ǥ��>��\c�[�Y����=��';hjh��ɘZ���V~��4k�-g�_G�=fW=���l!S����Lnm&l���7yp3JT�m��N�����<����Sq5�͎���zf����Z�	{j��F����jbI��"�É��T!�gi��+Ja,�~e9]��?L�^S������
��$W�����.��Z�O���]��6���N	��:a�Ƨ����� ���5�Ӣr�g��Ʌl�u��+��Wʶ���kd�D��1�ʺ���8+Tsz���-K5Ş�vd\�g�*l��p����ON�������_��Q}�;|�BX�S��',���8���z[Ϯ6�������W��bH�\hŷ���ǰ �M�����^Rdo��Gh:�z�)Z}��.7�Y*g��rI��:Q[�+�O N7ЊZ>�$�����J�c���~��$��A�D*,��6��'oam�k��6���#�2]�]f(��q�|Soԣ[���e}�F�cG�S'a�f}���[T��yU�gS�*~�S�vC�#v���W$`p�߱�Ra���(hа��D���Sq�YD߽-��J��cgq��*$�Ʋ��ab���~d%�6�q���R7Y�<}m���j�Tm��\�x�V��� &0"�"  �(�P���F5�<
[W���t�2�v�:GB���;�p�W��~@�Wy��ѱI���(��ܰ?θ!� A�D��ʾ��zM��`X(Nt��g��L���
/]$hB�.�tm�xN�?ᗆ���gÊ�H��U�1#ρ���X8�7�KFK���Z!�d��T�#�
���~ն.cB 4��G?[��9��8�C�.��n�8̱:' ���!k�JKaZ�������X�m��+����8?����+�J`���X��E"p"҈єո�q�lIv}f��3L�f��n:v�8�L���<n��U��wU�t�H�Ҙń�Z{��b!u(< �.�t�yFV���s
�Ʈ�UI3���¡�������Og�
.i�0<VRV�g�V��{�.W����a���`e�`��^��aD)�aV���=ȩe�U��Ӯb�D �@ ��=>U���*�˄J�O3h����	x�3BT�_�j�,M;U��7�SZ!�dix>��Cmh�Of=0݂�&y��zΥp�r=(	��ֱ�s&FOd����&=��@�˰w����U��5�2�me5?F܎��p���Ī�ro���~�Z�C{�Q�~�	��'����j����*��"(�Ԁ��I�yP� Jo�=)+����|��k�nZ����J���<H`1n�\�����1A���ЀѼ�D���p�����h��X����l� ��@�_��{�(X���X�D:0���*\������^�U� �\��Z�\�B��7�����Nam�tn����5�ء�����H�1MT��kp��������<5Zt��#�8�!�7Sa��2C&I���u�����K��(ɱ>;܁8��]�Țk���F�y��Qmn�D\�#�]�����H\��d��f|UU$�<��:(>C��h*�`v5�)أN!��7�}����q�e���X�BJ���p�27����|}*��,�0�Kٲ=�|�ڸ���o�m>DD=�O��.�dR���8<�J�'A�v���Փ����2��=88�l"+��&e�#���'|�]u� :��Z=%hm��<ϛx���̐��M��yQ�`-*O�֛<���fS[��24�C�༸����7q\��7 s3fsצG��X�
��A���2o�J�v+�Y�z�Ö���y�+w4���X9ƃ�"��p�.��|w�[�z7����4u��f�`>��f�)&�Q���4A�_�ԛ!S�<d���2>G>g:jݙG1yΚg&�{���F�}8�e�����u~8��?Y~��y-��)��Ç
����DN��1��$t��7p "�+���2������,�y4 �
¸6b�庆B�tN=}(i��bvU��AhR������uGm�q�+v�Fx�1pI+�И`������,yb��\�yĂ?��}C3��[�4�~�q��L�o�H-	&?R���q�mU2�Yӏ��Vud���@3u�����كX'� @��q�Z��D���`)R�����JG妀?g��t�-i��o���=s![B���"W�ޒ�Ѿ���TM��+�nӇ'q��{dQ��,>�/o�d%���%� tL�L�H��֬����u�:���c�P��i�v��p�������鎵�#��nH@�~�p�\���2�����h>�?�K!iL�L����9�	V�5����u�af0b�@&W)�1��(�9[/�捹A_�q���<�}>�j�G�R�@`��J7�' l���	"��;=��ƫ�rbW�=�"S�A2�j�u� ��SS��.�	�F����zJ���Q��9�Z�f���c�%��m�4�/�%K��j���=��T��5�$�Cv��B�59��� z,�KЦ�o
~]c��r2�4�4�O�n8��'��Ig�7h���5��>������ޛL1`�*�%qCc���{�7իCS�V��%�m)�"kS8M��Q%���,�� �g�t|��'dڿb�^<�&zBC"{��4�C��H�=���˫��A��-	ѓf���p}�c�ީ,�� �?�f��ab��P/��B��kܬ瓌��ʽ������e�!X#���lG�0�9n�S�����������,�dƝ��Ey���Dƿ�W�K�F�&��6zQ�D�8� �Ay���k �X��Q�/ �e%����Ԉ�BD��;�P��� ������6�L>�k���ȫ���@K�gdΚpVvk*��9�v��K�<!�GSއ�ǫ����(�Qf��* ��
���u�FB*�K�?�8_,�&+�p_�Z ����z���Io��\.�;FpK˿����'�Ô3 ���ǈxC��f���mD,'�N��|\�]-����L��������;��^����(�1	�r�tRL�P���o���,,M��R���Z�r�Gs&��$�����ͤ3��cX�N�ю�9P����rӰŨd�열����2u���[1��;�g4�h�Qy�;Mv\�B�$���f�y^'�<~o·5-����+�.�̟d���Zޛ���NE�F��֔F1}I���Z2�]�V���\o2�0�� tsă���TlV��k�g4�_\�dT�/%Dջd���45��F#�,x_��� w�]���!Uf��O�.�>S�2}�.'5�̥?��x�<��N�Ze��J��h�����  ��%20�Aj�P�+#֬zy�N^hzt�_�*�^�'>}j(�y��O��~'�L��ǩ�9�(��2IJ�M���7.C��<����C �kq�p����\W�|wW*G5{)�����5(�Y��e�_�N
��"4nd�7�=ˀ���-@��
68�׫�!z�����k/������ckn"m������5&�|f�J��B�������u��϶P��m�Ya4�q�F	�Gd/�ĺͭM��	͏r)�y�­$v����"p�<j�M��[���~̆�&��P$h���n*� ��9���/�� LI��Q$?�?���X�y�)	�<��T@?'R���=�����KV�	�2¬�ځ����ҽ�����.��)2LoE����g���bh�#�\��,��J]I���r�q���Y��
�3�F�n|�-EX=Qj�։�\��L���:�q�ZNx����E�����N������M0D7��Y���[$EFc6�0����8�f��!��0nA"�x�|�S�Zz؅җ��-G9 �K�Els�g�$U��t�ퟮy�J����{H(�9ic��8D����Y{�j�k���X���(ڰ���*ie �q�do(ⶼ_�_���s����k�+�/�(��R��s�?a�_>G��7��9L�=∌�t��������Qp-5sg�K+u�h�q��o(���Jx����_8�x�����va������
��r�[����p�b��!*�����+�l�H���og����1�l���Za� Ƿ}.�Ԕ.�,�C+E�AH��.���8�vC��౹X4@�"�a� �YBn2��J ����1p�����{�����l}
t�c��ʘ��8jW�C9���W��`�c1�S���L��?t;�Ѥ3A,������u��$��h�@M����%��VȐ��LA�K�h�s�UV�?n��m�bv�/������w��_�<UsHW�"��Cw�O�I�%�	�P�Rf��Q����j瘀���1�o���ۉ�R6jm}�)K�`�Z��6P�ކsl���/P�otU&1YS���H��0᠖�twȽ��a��F%RU���<G���G;�N�xҕRz���e�S�mt��`�V��	��;M����<�Q�E�G���w����]�g��͂�/(��f<���S�P���d'%�Nq9�?�����b��p�Tޑ��SLG��l��1���j��ħ�������=���Ε�ޥi~N[-��2���y�5���$O+qFf�CF�Z�J6;��>�~!�.|�vQB��#��g/
��v�p-���ǰ�����%��|�{ ��X}q
7��ɘ ������/�P�e����k���y���r�{�����	ԩlr�V�x���9���h�yY&��E�ia�]�iht�1~h��l.Ua��g0⺃n���~>53^/O�1o�n�uO��:o�e\��}g�����oS�j�8Q�L`�F���8��tt�34�cܐ~Ls��P���ne�'I���Ƨ`�
+u=��e*���h�(�p���]]���geIS��� �"��ϖ�,��)�����Ϭ���oYcIS���!|Q}���i��e��@+ܰc��:.�K�E��5G�Ob��C��绐�+|���Y�{wV.{�S�;Ռ�>q+��˚7�{�|1V��fBeX�I�}�h��:Ff��Y���Z�ɻ`W5QG�Z݃��nVBƥ��B�/���n�*g������n�]���L(W�J�Q��(b����7>Hv�*A��;��)HمN[��Ӝ��A�i�/� ,^��-�?e��Rl��D�R��.J=���?����p5�_2���؎���]��AD���P�PI�D*,�g���$��h��:�+c'M̒ړ����K�+hwf���i4Yѓ�|eD4廬������eK΂��G�B�ū:cj�@e�Ǆ#V*�0�]������>�v�~װ���U��Z 5Ԩa�&�HOJ?���fP�I�/
o��A�*ʉ�ƥ�{��||rA�'��QV��{�"N(iΊ�<���Y�h!���>�q��W�xcYb����*S4�NG����c��MY�6i:�� ��[V�w|DC"�F!�����������֢@Vac7a^�j�O���8PG�s/��kZ�Q����B]�S����q��w��%h��G��ݡ�x�чUs���o-�o�Z���X�i�)x�n�,�+z�����{�3�����hQ;���#�t����Z��y�I��]��a(��ΉW�	:1!�j?�����
#fൔ���p��B[ʪ���9�����Fl����s��u���+3��ݢ�X^��^�0o�ڭ�=���3��<1���UI��W	�����Ŗ$> ���v��B�-��tSʏg�Ѿ�?4�	�w;�*`�D�iJ2i~�]M��gH==@$x)Ri�fѦ�r-�Av�N
�:���"w����A�!ñ`�l�������yWU�V��{�8&�h6��w� �A�)��(¼y���d�)|hc:��\�!c�pO��I�'|�k�Po���*�|(G���Ɏό~k�P�JSQjm��<���"�o�?'����{qP���Q����3$i��l�.�}�8���5e��_�Ӡ�_L��L�6�*������(.X���Zg�$����ŹZB�x>���Z�&�A��ߕ�}u�^M=U�� �{~{�n�,:�4^Ɗ�?Ӧ8�0o@{�˿�;��f��/N�ǜ�%�M<��W?���%lƽ U	�����S���}34��5V�M���A�ѳ�Ł�+~D�'Y]l�F&m��ճ[-J�N�[C�p��&�h��w���Х��6VZ�	��wN�/N�R�T��7�DZ�+ё�&k�b�h$�����ޝ��mm��t��� ��UGe][(�/t�b��Vo����ݵDH�E���z�GLL�3�lC�����!1�r2U�u;����)}���"@b��>�\��E&Ma�1�AX��HK,��cպ�3���*0&���4�P6�L-���)\Ӵ�7S	^:5U�a��+��X�VnH�i�$��U�d!���x�2�!��'���ވ��F��@��z�3�ɷ��Fn���P"bl:1��߄6��b](��C�pl��̱6�«��H���ܮ��A�dY�&�����#�](��H�{����pǝ �5�U㕸eo��U�C�m������yq$h L��2�V�l�XZ! ��]�5���S��gb���J *�n|�����o3�����Y�ad�%n�@�oNfqu<+�7C̷s�H����]��C[�Y�&s�<��^�l��:5��H��3�~�{OJ[�������0)�jtf�Q9�|�,�y�����6빊z��7��_�+�'t�b�w��̜��B�c���xo�(��qM���]���x��=�-d@���B?��ѵ	�^�R��![�߯�w�Ha�̑�/�Y�5�;!��K��l��%]�IT�$��Q�	"�,��c]����������Rv������D�:��Ō@~�k6�]��X�*[2B��f��OGL�!�HA�ψ6��D��00����KW <�׭
���:�D�I�ơ��=��i�Փ'��,���R>�	]���� ���̏���u�R�AAFlzͼ`/���w`}I�xQ��:�k$�p�6�O]"�δ�w�s�� �ɾ���q��k�j����k�ET���K����@ɉ7�w^�Q�rq��"1�z����1�_��E��f��=��=��b�8��Y���{�R>��y�u���qұ��A���N�@*��Əv�K�++����D��Khޣ���H�0 �-W�'��SQ���Y���U�}�r�8n�c4���"��t�uko�8��Ʒ�6J����&ޘ�V�{W��
@=��ğ�rw�����t,u���C�}��F�ً�ɳ��梿�i��Ԧ3��P��u�?����F���F�즂ˆ
�P���An����ڗ�ű[��Ys�U�'7�а�I-�¢�>r��QQ*q��s��i~�6�n�m������S% 4��u1*rc�j ��q���s/L�U?a�̓�͒�0M� P
���F��<.r;����1�F���@�����e���N^�� [�k��\P�l�~�]&��э�|{�x{vީ'(H���6FssKP5����](��I4+T��'kf!��5&x^R��1�u�����T�t&��)u44
3d��ZȞ��M�����=�]:���'i��"Hb=S���|��D_����U.��/dLoD$˻�X7(�l�AF���"�.l�A�-,v�ݰ6�^��^��]��"�����F3�}=����f��-�h���^�x�cD�4�� \�����1oͺ�yg�&�A�&��
g9�a������> I�hC�K��E�r�ޑ���4�6��+���(m7����	
�c��E��ݶ���0�(1�K�x'p�^LQ0�L��b���3U��u��[�i%����/��f�	�ج��M��I.�Qѹ��@��?�-�XU�SX�a��j�IUr��KQ(��m{�Y"|L-&h�pmF�bn��5>�W�48N���c��)��zN�0;��]����6��
��yp��^8)=m�m_��3�':82��&�=�J]��9*�d���.�#\?����U-�"Vb�A;�t�M�9�k�&��8�
��v�5��.>��9e��s{�V�W��~]����(����(�ߦ]:1���/���Y{����8@���4�rV)�A��rݺ@�7��B��R� Ŧ�lz�9�=��o%�
IoN�ͱvORXϯq�;�w���S#��TN�䔍��Qw�M�(0o�
�@�!��-E�dכ	�r&��=����'��n�〝]��$��5��t�ΰ�A��(vlk�J�Ù���a�R����`��Ϳ)*t�Mp�|�FHQJ#A7M�ĺ_?�ls�����O�m�2������Ozn"�J&A.7��-�`::��Zrfw[�Jzt<B����0�����W��X���`w���j{hy�o�"˨ �����o&��ك��
���R�=m�#��P����`��ٺ�w,C�K��Ǻ:���tܣ�8���$���L�]3%�>�f.�2m��y���3,����;�އ��+v`�"����;��ٺ\,��mʥz���ވ�� �>�dP	���o���n��v ���֑�������&Ahm6#��^�R����w�S�l��>�dd,������̦
��B2��sg�opؚ��`j|ڹ$!���I�����0���?�*��j�/�v{�XR���Q>�*sy�Y�8��c��ރ�ە�|Á:K���7@���*�u�Jm���a���	[�����*~�`�O��s��bX���R���G�������K�,����ӡ�x��ޮF����n��������#��QΒ߃��CӦy��c��bߌ��y��w?jq��J�f*/���̢��7�]�[B���H�/�%��/��[[K��`��8鸰�?���5+Z�ȗ\?�
���N|��"Tx:<7S���0�s&�����'����њ&Y|���s-��)2k�PM���R�qh�
5>���GʆV�$~��A�`����!�}�&<\	��s�!?m)� �?��T�w��$��(��t��b�5+�y$�O'=H���U%
��)bc�Fm�7�����H�,5�Ҍ�/~>���k�r�k��Rg2>�x<�Ix�];�ɿ��>�G�4�l�KUi9q�5u���=-�E�ʬ�v�@n7��5`�75�Æ��`AԌ�Q�
3L�w��*v`�I�f����e|͘�Pv\�<�������)3�6�^.���7ؒ/?=�6�Q3��=���e����X �ծ��d�AGbH�N��	�����x��(��K~K@���T���(}� ��hZQ?hb7��D,w���l�[���d�X8(3oܭ2��ȇ� �`��Z\�^f�oi[S��n�`ɧd��k�j|��ɍ�VZ�S��0���=g�G1B�W�\��X_��p�ت�cӵ)k��Z!<5�{��S�J:c�]���_<���R6z�g�	����e"��� �<��˰������.�44&�#[$$0��b�����?٫���J�B�ʤ39�̔s���!L']k0�)K�O$��6T�1��n#�s��b/ ��G�'��HD���Et�G�Z��g��I�$����s��xo�&��P?�#�5���t�$��W��=qUU��q�%�?�s x�Ŷ�w_ O�����~�cD��9`��vG����-{w���)h����j�}#�����F����68o�3s�Տ���V붻37��[�?�.>�ۡ:R��,�͹C�0x���٦&�"h�vOA{��*y��C����%.�����O��[���|�G��E�\���x #���f���l����Z\���P+>���|���G?\4�X��' h�Ym�������)zq����l��㱧����ɪ�p���?3�S���2+��ڛ"yJ���-l�}Y�v_aU�5�����R���* ��Gr;|��Ͼ茄N����5䧡U�l��?q;������"O�EEx$�Z�q�WW@�bl�FN��o5�OQ;aR���R���X#NU!���ޞ����]S՚�%��p������nw��s�u��b����7jN��*�6*Fv�P�s�D�{H�m����aI��m�~"&�����|s~5�R�W�ɴ�� "\#l�#'@.�͆�	@-������������h\n�:���q�\P��Tn&���O���m@��sW�͈���lR�	v��p����V�u�3�ʯ�#���0W�ˆ>u�T�b���;X�)���e��)���cJ3x�'F[RB�K�G�J��q���
2g	��]�g2v�k80OH�_�ϢF~Ye> �*Ǳ�k�9Z<Lǉk_�h��x������a�{p�+'�2�:~:H��A��b��is�Wl�[����|K�v0C)��,�ɩ��(��߮�DY'}9Mxr��m�� ��:���9z}�&Љ���0`�K���6��(�Z���?�d*��~Nu�U�����%V�-<_;�<���K�|��!D�����L�su�⏒��ZFg2��o�t�#� F� [�I-�pq#�)o����m��Q�5]e=Yf��V.~{
�6+�ܙ��-�=ԡk�<Hk���&�$je��TP�9=u��p�`o	 D_��.�D㻪tAinX�'���{�rt0<�ܘEg��xǹ���l�\_3G�������_Dȵ�&Ïs(���8'e3!��:����P�>�R��&�Y���l��l�ީn:���@iҋ��݊R��M�~*�Ne�&r'��� ��_��ؾ���:{_aP���9����K�Qs,J��"���w��;f��X��y!u�8Il*�OyXǑ��@I%�K��'2��>=�T�����ʢ籒���	,nY���d^���h<3A� ��HW���h{@Է�>]V��ܹ��,�%�E��Y�*�� _(u��a��9m2*E�!/�R8:���l��8\3A|

2va'0�[��3&��-.LƎ�I6�'W���� ���1�+7�`q1A�^�PH��=�� �n�7�N�s.����5_9�@$�t��:�WW\��*��x�cW>�JH��r��'G0�_�K�X�,\2����{����&tE�oJ/����vME_���B˚���o$ʗ�����/n?�������8־�u6G��R�tO����5��s�/ɐU����`�ʎJm44RՈS�:�#?N����iXhq����ͫ��8C�v�R�}�\�ř�X+xC��~O��_��.�����O��*��|rl��&Mc�46u����t��0~��s�8{F�t�x�$��gG؟��'�&�+�[������%�ڦ��DP�j|Q��ao3�b��6�0hF]P�P��k �xU��o���d��ã������+/�����W��� ��2Q��B�R\���K�Gm��69�E^p�.�u�a�+rs�ls�˻4��(8���Y�U6��H@)���]�C�4�~"['��'@��f9Μ*n%��A^�0�G��jR�����v�J@o9(��o�;`���I;G5���+g
�����m�`�ޖ�fO9��J�=�%����pӦ2�SI-+O�AŻ7���ʴS��xj<���/̥�f�=�E�H���A�1���6�����s��.b/�BHf�mx�����?n�
ܢ]-���[����b&`���$�E��eWl����'��g]�h���ts
KP��C0q���߰RF�M��'��.*.r����A���BJ�	 X�� ��,�	�ck�3���%�%n�[�NF��̵{+��Y]�	�;F7�l+2���((�*xUd.V|/�E�q��,���{�ė�^����T,_�#���N��7�(<�CS��b��8�E7�j��p �l��d,�����۷K5���7[��������$��o ���d2�����d����ޗ�����v��xi��
{2_�s�8�� �&��A�YS*�~a�e]� ���v.v���V��\b=����g574�E!+�6��­1<B��>��⭭��vu������.��ɺ1ҟ�+��Bx�*.�����]�h�<�'�V�{�!�I��e���;/9h��r���ͨƂ�{��� �Fc0����Ԣ/q�vw���'n��U�o�MI�@��n�F��Y,^1i�
V�z}zvH�[x�c�A��y�}Ϙ��bM���Pe��������ehsw�p�[�ɕ<��=锔��M`L�#���_����]eȗo��^LE�� Jz�#D��o�9�u�����n�����ph]��A��
�iDK-���yނ�%�xW����+�t��\z����caZE�����m\�<��P?���^g�"��Z��-j��ÏyVn峹��?�9��A�la�����'�@�6p�S�M��c|��X0��̭�A��ՂN)��u*��rʼlo��˰������v��i�n
���?���hW�o�.s9�s/�Fd�ޭ��P�;3w�������t�E~�r~"I�ҫ	��7��D�F-[�{꼰'��t>�G�-��2�����b�C��/ '��@zb��Z4�r; ��/>�G��*��!S�_��}�sAaj�����9��?/����9��$�OtTi�O���0�~vV:
�:\*i%�5����iy�I�:2+:ו!��vAM�MW9A���[3�����(	�0�4�d�;�cF��P����!SM�pzd���߷~������4M_�F�+s�"hoq!W-���a��vFW':�HU6�Lrg,:��(���v�j�_�b�i�Nq5����D�u�;���}#*K�w5->mW_W��'�[�r��õI{Ӕ�f����Z=�8ȗ����y�S����)��X1|Z�.�`�t��Av')����G�!�d���A^݂�pX8�t7��5AC#��)L��1�H9"/��wri-�{u�����
�7��� U�� %
�^����}���Cj`l|�K��B��! �`��_Z`�W�C�����`�L�l��I݌{L�#�&�nD���
�x��?��Q��$�I�?�h0#�D�EZ��=o�ܸ��uUnOp4��8�9�*�r����ˑ��1���L'�-8y���o�3�=܈Uq�hl�W&��d�a�p5�u�RnK��zC�4�d*돍�%�����]��޸`�Zt��-j�z�5���YPXV�T!>�8��,��:O���8����Ж��j-Z���v4"�ܫ�H'��vV�.�qy-%4;^��a~d���t$� R�Q2���[��O����P�^�����ς��Iۚ-K7��?V����0��D���t>��>QՌ��������?�c��!<#[D��Q�^4N��,݋=4v��mm��&�c�RKL�G�xr
�Dʐ��i�ύ�_Y��[0+��� �ދU����rB�wc1`b|u=U\Y��ć���[DGO��[o�mh���C}�r��o3'�&}~��K���8�A�܀;�ǩ`��e��9%ऎ�Q�5�Y������\�E�T����z�����M/�[�cBj��m �Wt�Gw]Vu�LS��>�F��L����2���-|�Hj[�,c�G��\�&�4�{�2���H ����������L�HU�X=�=.�B޸����F��h��z��+���jK���jbf��|��ܕ&�}f�y�h*yz��A�s�G���
?x$�~���l�|�3&X�	_�7h��W��3s�;A��F��iL0/���+��	o���j[#�WW:N.MB�:;a�prw��!b���<z�AM�������Ǻ;��),N�a�����ޢ�A��[�ݿ�ԋ��#fx&����1ee{�m�t>�:k���0�]O�������=�xga���)Jy/�6�~�urm���8���'!��B���Ty4����6�ա�^�R�#���	�Z�A�����-��rv�-F�Q��,��<�׆[>��;����́&f5�����j�WVܸ�$#Kf��Y���$�Or���yX��^�<�F�l~4f������d��'q�����U]�g�W�-���*�f�*UJ���䩢lǷ��t��Y�t���΀y����鱋7M�4��T���K��U���H�5^�=(Ŷ��~#�X�L��`/����P	��bS�յ��僘g���J�������MNq�����[U�$vH���>s��gx�>GBY�-�pӥ�?����*��@�	�Š6k��
����5u5'�g�=��g�ʦ��� ����hA7���������–�1V��f�'Y����.���M�4y��n<�e���_6��[؁�
7ބ$J=N=��Ԋ�>��4��@X#������ȱ� �#>��5��U�.���+11���ͺ�@/*��>�m�N��*I��D䧊�FZ��y��c*��Ҽ�&�3'�[c n�N@�[0�Ӹa�9}�i�
�]W�@LQ�{��$�ͧa*���̶y/�R���bǍI�+Q�����1�#���@M�X,}������~��6z[�L���E��BJy�x�ǭM�X4�6����Y�p�>��}�iagQ1͒��,�j�U�~�����i�`��o�a&sBλ�f/b'Ѐ�'n�L��<k~cc���ج��Wv\��~��'�*��=����}	?�C���_LY)pjz�i��t#v@��E��)S�����j���zI�Q�>9����g)���w�.E�H�r���w	>�n�ɹfd_:���)�e�G����uf�K��Fu���ݨ>K+��|��h��!�,�Jt�	�=�k6,7��b1�>��~��z�pu74BAl��XF��)2��2a�����f���H�P���T���"�K�I$�:R��sL�!�D�����$�tK�֛٬#��U����z��7d��R��g��K��0;$IP��Rdw�Ҷ˒/k�إ	�N=�:ʾo�spZx��S.�p�E��ԋ�ն��g�H�B�vi���](�S����6�ֳ��t�a�����|ʢ��<�5o���O������
yw��ٿ������;��n%"P��>�GnoO�ֺ|S��O�`1`�(�rc����иx�V�+E��6#W���� {�����'�z7c�ӭ2�[B%x{�o�2�Y�v�����zV2�H�a�f@��E#����Oi8;�'p<���x��XiU<qW ���!�Hs��Q?�����Vٽ�93!~MzH/�<KH�dr��J�:=�4R��ԓ14��D��gu�-�i��<N���i�c0y�
�0�����k<����Xe-��U?M(�
-�c�:�e�B4�YOM�Ӣ�4d�6���w	����X�wT=x\>iP���	heSA兔c)>�D%P@��4A�μ7�2f���d���DEm�]S�h�Ԯn�=�S�������9<�.�^�z��(H�
�������J]\G�cx���ooJM��s�!��j�BA9�ǥ�_�	:�4�cB��j�.~)G��JCf�h��+^�2�7{��.Xp���z�������8���P�89���d�ApwA�����e?Ն���G���`�4Q=�	�~�y�T�h�[�
��?XTYК�]M�$�F�o�*68���K>�$���~��JC:E�������.S�q�� W#�!T�B�8��>��I@FA����dg��ƹ�$�I*��>��r����ѬT�;Q�(�E��P��!<f��
���w͘��@6�Yl|P��4�6^��Dkj�cNb�����(�i���Z�q����C�Or���2�`�8Ap�b#X��ٷP�����b�&1�Ei�uS�c���m��iGX�vC���������d�20�<L��%{k0�����<hb�)"F��+R�������	5��ڸ�;��y�=J��wγ�/�����z�s�ρ�	���5�Om�C$&2��E�9�G��" ��Xcb�TF�h_Ms�F#�A??*��e�ǖ�ۊ�o
��`��le%�b�=bA���?�[yT��M�v��G��<C�
�����s^u��ra?�(:��@�J��dv4y�1�i�k�/�k���JZ<\eJ�MT`�������A4���/�xz�	�-C2%�����F�XqȦ.������g�0W#k���K$����Ӆ*��.~r�9+�\{���?�����5�ZT�1�}9�D�H�yp)jN8�����okLIG���{,���~m��!`�N�g����ʺe�+�AH4�7]y���$����/r>��F�'I_t1�WT����>/�+W/��9�pՖ�--�Fm�3���ڸ0:a�+rd��x��d�p��K�)�'�Uzm'{k�A��1��{����N*Q-����2
�_���jy	/ߺ��I�
��rh���̻
�
+�װ��u/Z��,�fע,_�IF+��{�sn�l�ўCD�O����)P~�X(2qD��z����c���{e�̗�����u�_y^d�:Y82�0�DL@~c��������.��)���{ANe9J�s�)�Bc�}I:�JVa��m$	��&�)2�
�Be��!�r�B�y���d��hF�Ӊ�2`�6�i!��I��bQ~��pj�`*�^ޡ��st�%[��f铙=�C;�;������8vS����$�K��oJ�,�m��ҬR���η�a�6�e?�]�/�Q�4yg��;��WEֿi���}.�s��18�[���������f'�2������>�����f�-5�iK� ���O�i��vpZ�X/�������:H���IӭWK��YQ��?It�n-�Z�1�D��E ���]oD�`G��|�W��H��yq��b�`��=���,#�6x�\��X��}sV^�H��$O���	b�
F�}�1����R���\Y��qHW�԰7���k���Z���\=���v������@o����Z��^@�G	�T�S�?@_		� �~c+�:�n"�O�U����;d	v���1��RPӕb�Ԃ7�Qa�:_C���ϧl��X�7NMa&a��}��R$Îm��<\'��$����iK�c�-"�9�U���ܮ��;��h��|laɱ��$������^ک���)�V�߮g����>1R������9�-�$�c��tg�4vp�Q�.�r��S_�8�Ѩ_5���I�h��Ѳ2L�j;<��W:Jtb�vG���P�>� ������~��'��t�y�a&
���hn����Y�P`���v3��4��[g�)z�F�Q#�_ؚ�&����{A�Ł��U�z+��� �X�J�`��N%���:�!!�d3D��-8L�}���&1t����s����y��W���>�N d�P-l ^��;s���o�i�hN߈��8�?��X����Ͽ�m�bU�b<F(&�˜���hI�{,�!{Ļg|���X��WW=�+1�#��WPV�xĜܰ)�0��I�nc�����[�3���P׶&���7���T��w�~�|��%jM�Ql��\�O0'��B.�ڏ9����N�@�:�Ҕ)+N8�6�.�x�V_�$Lۢd�W9у���N_3�ׁ/�p���k�W����\�~!�+�I,ʴ�w�],`��%��r��잤�3�vgBG$���s~�[[|.��W;��ulg��Pc6��<Fg� ���8�� #n�x�g|+D��f�Sƴ��/x��n�]k ��������u\d���1N�)�S��u�S��f�M	�ï�G���p�j������v��Ց�3B_}�k1@,�:R�]B4�g�G*"�v���ԑ���=t-
{�J�����SD�`�e�����P�HO5�����o�d�ƹ�Ś�M��9��ޗs*͏���N�� �9%��ka�m�À��nv[oD_�>�65���+���L�^�\�����P���l��9�E��&P�6A�?K\'-�졝��c4d3�3�!�{V�l׶���n�s�e3��!;LܲМXq|fS�u�( �@���}�����L�P�5N���Dv����5#��tȆ��������5@�j���!w���󸯷4�)!�F}@��cO���B ��nY�k����7�AD���C��Lz3ڗ��w^o樻d,��1y폣ΛؗK6([����޲������:j���`|�eٴڳ`Ν��|]��8v �X�����j/��;��6��y�>Sp�"R���nk']Z�������~[����!�sy~��f|�OR�3B�n����M�n�����g��SՍ� ��4e,c��� ld�w�ƖV��,� =|6�O{� S`�6n��mu���g��KIz���^[1X��o&\e� )��j|�gU�^��I�?�A"%ڣ8�l�-vYD;Y�}�zŝ���<��mJ�1�(�/o�aZGk�"�������;}�O��V=xM�갂I�e2U�¦�Uy��d#o�O��w�0;����[hh��i��اb���$�Vز�?�)��JK���s�sgG����5�kYY|���fM��R�VRQO��?9�<ra �[����=�p=�t���Y�ٞR�J�q��XP��A�D��]��X�0�N����'��ly�#pzIRh�y����lz'�w����,'�:�Ur�ǣ�m"Ʒ��=�;�\��\�rU���2��Cɂ���0��Or���g�����Ъ�F��J;gP�
�_N1]z>�Xu˕f��|�&J�X�V@��:����N��[T��N�x�Դ��3�x�2s���y�a/2C>��|8̎��J�7����`�>c�~ 坽���oZ8��S�*�"��b���A/�Y�(��]J��{wn��a��~:܀4�A����R�5��̽�W5�fk5/���,���׃[���y�+�'2����}��@��:���9O�����h_�K�s�����Yo�I���+}��.Iw�SE-��b^���%W��:z�,�ZV�&�f���Z��oK�L80R�t�`���yYߩ�SXy�mG��hR��Q�|��&g"�o� �ݖ�/=eT]y���'m,x��m���g��.V���#��D>�@�{�rq�x��o�yV6v��K�(�(��a��Q}*?X�<��Moz�
�m�W ����Z�=R�IɈ��־�c�)uH0��k���-�4�ֈ���÷e�k
��y���5�ɂ��3K��D�".	F�L!�%Pzc͟���� �Gc�%�{�ld��� �o�~��}P�z>�xܫ$����ݟ<>�Kwx��ǘbz�r�#4�)%V���=E�����M��OY%���������������~�O�"2� 5�j���t��ҡ�o�g������v��i9@{��#M�@,,Zh�v��!U�v���~�s	�y! ��\��r�6$�p�@���@y����M���Ud/�!�c�����p��b:	�-��P���)	<,R�7�v�����=H��tp�ծ�ab���{����t/�˄�,{k��n%w{S�|���0�;���>�I�^���!n"I�t)��-�[�D[���ŃV�����3t`KQƫb��P�����](���B�� ����(������On�w�8:o�'�Y`�v�w��YXd�|y�Y��yNA!�^���6����%���m�)Z�C]D���X��'��7�N}�Zd�	v�TE
>F�U����il��Uf�,�rYN�%�"_Uc����b>ȫ�9*K���$�4�RηU��]a��#,�����֓�	�i����@�;ATW������mx-i35�j�3����Ai�ӳ��X�����L�����!uvb�����J��7�C��<�2��Iڈ	�a�⬠��L��?�G`hL%c%�:����Z�T��#�������?��a|�|>�Q��� �T��V1wEk7�H��J(>q�Z��ԗu��ڇ��;7{q�";��1���^�J���Y��s�mm�(g��RYjs�գB� ��NL���a�`�6�J��"�m@����߼j���{��a��
UlSd�	ngG75�G�{Z��߉����
o�&D7=��6W��#x�ILVu6��M�;x"�_rf��  �)��o�2�r�㜩ɜ���?!�>�,e�T)(��G@_��k��ͫ�c"�i����+���9�l�|��< ������>�r=�Ȣ[�`w��
�F�~�yO�B�j�}L���u�oڨ��?$:����{C�u�=�
&�c�������uV�;ݬ�*��H�KZy����?�^�r#H�)-@}����E�k`G�� ܨ_Y�uo�{�96?2A�3+'��������S�m[LB�p�"���5"rL��v�A�εS� Dk�*��s�}��;�H�iV�����^^j�z(ik���wH�^%|��5�ןt��Du�\���f�����D<c�$J+<;�{jnڋ���*�7�2M�14��¡��+(����y���{�A����F��Z #W��GŢ��F�M�SCO!�FC�e��sB��1wSՐTCF�p�&H��[�����Ù�&��}�Y�!��j�2�& ��7�I���/��d�=�p�����n��b���. �w(Cd䰽��mPLIG���=`7��r�Γ��P{�eZO9Q�q��6�x�]"I1*x3@��X�!��ӺЄ$���f|w(�U9��������K�|j�E���B����� w��Q�j�)٪�������5��T�QV@��<F�C᭩�C��z�0PWES�59Ą@��6o�i.0�W+1�J��}�[�
�CS�,�_�1�QdD{��Vy�믚�*�
t �V��2�5�G��o�u��d�=7a�����R5�_z��qCe.^"���7�G��pWQ�;Z�:�]C�Eݰ�R�>��i�����&s��ʩ;�,Qm�]bƪ�����ύ�AV����+f��ԑE����9q'��]�P+����ͬ��W�"�x�	
ꤋ��.@SF������VU��R�����]��2-�����0�E@/anR �lHtA�"��� �Y���A�ʃl���� 	�Z��"��!#�q~�]��Y+c�y�C�}�0ے���.���~mJ�HkA�^o5i��_Ѳ_��(�d^�J�C��U��R�Gk�gc��s�"T�!j��?~��.Q�Ak���y{�[2]tn�7K��n|�B���e�eY2���rB3r�Ƨ��ᒘ��T�/ֺ(hܝ����[F%m1����'`ZV������ٌ�z����	���t��_v�:8hY�g�R��w����Xx��X��ܬ�W�h�-M�a{Ne�ބ���e�GWYڒ?z�q�W�_J�Gj�uDĥ�*�c��ué+�O���7xT��x�1<��`_�Y?��e觴���0��e��9f�k�g9x@7uN�h-.#��~:7�2ڍ %�,�Z�b����g�q��L�{E�����r�E��pS�2Y�rD�������R+|c�ȁa�/7�����,���dS��g^r%@��1���U�)[���%;M:]v�& ��KAժ�ǽ���q�-*D�ʰ�Z��o�؍n�!	��.�0
m�������9���CŤ_�4�I
�k6��U���:��>!�4��T\䄐 )^2}L=�M�˴��0 �0�a��:����"�W���gTE[0�.�%>E�˕i�Lo�h�S��O��S6���T*S��4Tt��5Ln�i�y���o�-s\Y��۴��3���Zm��!��*U�oG F�!�}��w���C
߼���7�S��R.����+��m��&��@	�a�VÈs�Ţ��Đ��;�)5V}�$�´���[�\��Sn�2�'{�@��G945.�S3U��C�3�Okʛ6�.�6�l>�&F���ړ����KxՃę�q��B�5L�!STJ{����VKs��Y�Ķ�D�����#G�#��#�y���B��dC�cIo0�`��"�䦈OO�$$�_���:Y�,���]�}x�0b���2e�a�<-:8���b���v/�&U�%YkrA�+b�1�)vu��Ef��>����ۆiTu���?� �s�M�b�jeZ'e�?U��!.}�
��xP���f��ֵ������?�Gj���ky�����n��J��Q�2�X��@}�.�z��	��:�r$־�ŭrv���Ӡ�t�`2�_��PI͑����<^��O4쏉�g�R�yrZ�v���}k��Kw�����|,��ջ(�I3b�C�Ra���,$�$��xC�@�x<����V����u�d��K)O� �޳"�$�5�V��Q��P}�h�?�yG0`�l���	%��n��vcU���Cm� ԧ^��%`E�̇ha>��a[6ל:�B�8{Ɇ�����)ں�
����g�`,��"�|B����$�����~�y��p�� ���e~��'� ா�lB
�I>���x�=�E�'�k���%.Kܱ�A[s�Mل�g^�q/��fD<��E<���ζO/kS�5~�����-C��O�n��(���p>28q��X�Ww;����G���fX���J,w�w�z`u�l�8.C���KPUg����	:TF�+8�7�w)Q��a<]",IP{qm|��t;�r����~��kf���|,�!�&st�zD=��OrrKYr�cҸ��>\���ѭ]2�8���3|�;�I�v$ �|}"�K�i�.��+zDJ>4�t0��>���#����9�Y
p��6?��{�v/诽s�\���kAg��o���s(��ke�6#��I�1�����&6��~��~��$��Q���$�'�u���0��;���#dǯ�%3�a/R~�5j��y!�P����ȌB�"�x�.���,?Bt����� S�x��9F�q��&��I(�����ݎ	\��Y��v#�̈́[��*��j�T����1��#@��=�`�=����OR)��K��.�m<[�u!��΅�1V>ڤUڐ!	�(u�؈D�5�J�)a���V�?㠯���s�nn����7��?���.8rs�xh��0�-�_��^a+�c1�5#��Q�&�d�Y��>Zv� ����ʺ�Zj#�HY~����ד����O���򿜫Y�󞞼D�/��EX�䦼.���7���Z�u}��&h��{�U��=�A�}4��i���KGA�B�?�Q�pc����²����K �g7� 6)���ꔢ�\�v�}�BI�ō���K�5k�<4�f�����.�i�tϼ�NO����κ��zt�u?��;��Y3�f�6"��\���Q���H�0ŮRji<��Eg�>CL]�A}8ّ��|2��ހC��t�㍽S"۫Iֺ���i��.��4U��8��MNI��]����-���,Ā��ϑ��.�P'��	��m�X�:�q�E@#t�ՅU�I�bSt�ﲸ��>�Qp�h��q��
}���2@��<�#y��:����3�cs	< ����CT�Yi�	�r��9������FH�/�� |�����V�={w��oڳW)�(U���=,Y\�8�-|��.��N��������b�l>�~j�N���m�yP����Ȇ:y>i17bS��q�żL��v�<*��;���V�m�j���*xʐ;��z�/Xє�z+/M�0
�<�L#��s�j]}��X�'�����F�g�t�e�x_�J晃t��S�r��?��wHa�U&�j���1������pU��m!�0�P AI�
�Oz@�0`/Lф�[ڃct�4�z�G�f� Z��oY�-��O�\�Ͼ�r	4h��ԹB�|y�*�L`#}
�m�l#ʼ`�ޱ ,'ް]d�,��%"��kd���.����$�[@^W�.�z�A����^�����f�_�n�o����v�y���Ŵ�ǣ����;�G ����i|�Ghi�b��V��ֲ����:L���-���0�J��F �8A�\Ң�{��"��.����ow�mw��?�ʇ���g	S �6U��i�;8%-_f*xL��O��2T/�]g����.Go��%[�@���m�$�ث(����<.��%�Q���90K�T{�Y���U�@��ɳ�;Q�d�Am�b�}�/�<Do6��b�y�L�kG��*^u�lG*ɯE�e��D��i���!3�e,�J7"�������h���)��E@���p�v�ݮ�$�>��NG��A�n0�0�S�� �3ͭ-+t�K,Ň���Z��>9'K�	:�t����e>���ǟ�~��X�>|M��2.�F��"9��ؼsC�Ɍ77F�q��Tg	�� ��p�3�p�y�;Jz�%�w��iova:��U�^�h�/�*����ie|ԬwG��J����#��a\��?0��w� W�� `\b�(�y4��&�n-T�tm��=�%n'�__ؚh��	�bĜ[`���L�f���6�L{���G�H�OHOH�������YJ���� @""��2ќ	G�C�%E����0
��ML��WF�vz�#&l��ns�Z���ͬ�<d��d=~:�)�_0o����)%����q�(���BÛV��㨬_�0�;nb���A9h�@���Ğ2�}��]�{��C�M�~MH�)�ui<ǅ]�5��^;n��0��Ct��.2R�8��?N1y�!�
z����o#���Zgd�D�1W~6@� A  �A��X� S�Vd^�r;y� ����zQ}��͢���J5�^(G��(��G�S$���Q���K��ңū<�0}���d��^�G�i���>�Ԛ�9'�+��Bέ��0�=��L��k�5��DIx�p'�U�׉�(w��
� p�/ڃ7���w��wt�4[5t��\�k�������e|���0u
�
�a=��٠�15���[���E�8l�x�4<v~HG��Ic�?����v�Qz�ז���I�1,�����^��3�E�a�Y,]63��z���uGH���sX�������� ���t�A/��1�G&�fT��Y#�9��i=V;��l�8lH��2P���ʻ�&Ţc��_ĖZ�ݘ���2d
�J�����R��MD�J��{�o������W*�[\Λ
�,�x��%����n���8���D�P�-�Y�]��>[� �ZR����b2��{���F�c�4��{Wʞ�r�|��rϕҠ*aԧ����",�f�3����
/'��_ÚP��Qy��}}QV� q�J���i�&�tذ���γ,��:<�<WUVAF��}=\D�fk�X�ۋ/�w8CO��9��,����+�`AF.�D��(�^_qE����S�hc���(Eq�7��d�FW[�Y{d8��R�x;��.�z2L�[�Z�KБÝ@�	��");f8�,m���G�g�5%�6�n���T���bF����P�7�jZ��m�r��+�������Aڎ��[J]A��~L�h�>�h�%iu÷N�u��?�N�-�Z��w�͵Uq��|~Y{M��Co�����9|�W���"��##�=�Z!4h�9�R+��M���8nе���ZG�6o��"kU�<a�BPW��:��-8�ࡕ�J`����7�%��F��i��\A�������+{*�a�~�*8������I��A%s���{K�m��_���MrV��J�����l�T5�'����y�p���O�����<z> �tA��)X�9�Z�QH��x'�����P"L�oeE
�D#��F����]-��y9���D���,E  $�$��x?�'`�`)��<�Ɔ��Z�֒t�K�����5	`�����rն=r4\���8�k᠊��k˦Ѻ����z�[,��U�[w9����f�\����A �ݓ� `�!rݫ�u�s�>^ǰ��VP���H���טC���gt�ن��(-��:��lRf+�S�_��C��4R�a������Z�K���/��ɞZ'c�����\s��7ж��M��_��C+��9��%Լ����������˒{��������^������3RWfX68g^uz�9�Tu]��t^�F��� �͊��y���k�R�Y=�PB���$Ϸu�{��:N�E_-&О�PICp�1�C"�ر��ّ�@�� k ��A3�N?����o�L��~�;^������kT"��7���^D�'A�@/���*A�߅O�8�4�A\�k�t�%�a)�ei-\��b�5�m����\\j(��-���x�Ii,6�d
�D(>��� )c!��,aַ��s�;�éz���7��K�s��*��"o�B���!��q$2!�8u�#-x��l?��
�����<��=�-��m�8����!K��ڑŕ/���>Z���@�f��G$v�m��A�� z�[o�F��96�ŵ�DF��Li�i�ڏ����bC�nȗ�pN�>-�=��d�&΅l3��␾E2�k��4����4��f�^�s�����(����:h��D.uQ���u��{�F
�pU�S|`����R�)vn͝����s��pWw-��7�Ķ�R�{y��~,M��g�����Ċ(m�м: |�����68���(ZP_��"��ӿ�6���/i�X��C�c���АK�i	���z~/sT�X�u����"��W�v=�$V�+B�w�Ρ�L=�,p~:n�.�a۸�yr�[H6"��͐�OD~�#>�I�2]��V��RZ�o#y"k�E��d{�:�I�UW}�`i�v��v;�����$��߫���.=M����-��{-k?b�Y۳�Y����s��dಥ��e�]@��Dh����4Nvto�^_=2fg���H
�S kO����!YX��<����Wp͔�Bj�i�4�77����s?��Cܡ8�|��� �e����;����Mf誴'��?Q6:�>���Cu#i�E�۰�fj��d�-�@��l��m2�|n�5�9oʥ7\�:7��
NC�@���u��֤����ӯ�L���2���}J��@�]K�*�Pc�̀����m�DE��~�E�σ_)�b|����=�Vbq��낰�C�J���yIfQ�׽X�X3@��PNd�Ӑ.Z5�'�j�-,�L��j9
g����֎P+�C)֖e7:-��
���i���d�
-ؑ�q'a��ߘ �)1�s�P�og:�{�O�"9�K�'��G]X|i�_��p�*�9%=%�D� t��C"���3�	��4�Y�����a�9ߔ���!��e����ItWl�I_�7u��^2Aw�hW�A
u�T+�̨Ki������%�A<ĮB]�b�c�x��qy�5���
�+/@��xbq<$�
W��HS�/������0�8��%T �H�&��e��Œs=��ܶ�kL� �y4? l3�hׂ����x���g�i�|:�`r|I:����j��:w���59����� N���S��-�&��������⋇�R�烓�J���� ��t�/0݋[����:�Dϖ�0L�Y"�H��Гd�C
���K�!�Fe�5�=׽q��7�C4W{~o�/a1U��kH(��2�,Ơ�b��iZ3�k�u L� r�3��i� s��5EN� pD܁ϷZ1x�YR�..-�5*6��ߛcQ�5R�(�"*@6��}��K���f�G����Oڇ3�K��#�+�&�P�U��vg;��Q�E5j�\�V�^���ߌ���ӷ7��u�Ni��4�L*P�Ȟ!�����ނ�9^��⢹��k��S:���n3!��@��R�^�����3D��P���@���U�yk�ĲU4�Hf�a�5�',��lX�l�/�@���dm4���9�_��`����:�R�nl��*�ܦ�rz(7�Ж�z�L��7�Xo��@�YbV�祖m��k	a���3PZ}�=�"(�.p˞L��te�[���G����m�WN6!W�~~�e ����Z�j�d���e�l�)���&�:�4(pFά�j�)^�4H�
���Z�ʖ���"Ǐ�d��@k?�U ��2��Ɖ/���	d[�
��NR�K��ϸc$����wr��s���O�畱�xf�"���7����/@��l� �0T6Z�ױ��� A���_G 1] �$y��d��WIs��a��7��SfvH�Jj9L�W��D�)��6�,��ZJVCy�>&8<���T3ǭ���3@�F	q҆(��uo%쩮��^F����&���K��]_��F	��aT�:xcA�'�g+a�|r�$t�c��a���ɬ�����4rU�#ej�Z
�.��{]�oOE��xa�t���nXo�w_�y;2H��=���!� ��D������]�
4)>�j5So�H86|�q�5���=�,�R��I��৙c�(�,f�m��sr\vb��bIaB��	vz���5ܧă�%ί�IUs��Xj%�N�"<�^��
I�!���a�j:��r(�hҭXf���#'V�C^���<�2�b�(�e=�v#��3f�;e���LƥfW�ķk���鳄D1��n��s�	�83j�]<U�8a�BYe=N��("�L�܃����*~ ���H#�z�{B�B��R�s����&��DL[�*w{&�H�Q�t�]S��ڣ�^_�o_�k?\4�u��86�^��v2*"?G��yYy�	�w�	A��l(5A^x�5�Ӎ�iR�z�K	��e���
�=DWJGg)_a7+���t�8}�� ���&����H2=�a��.�,��KV�/i5(R1� ˓�#"�1)W�;���b>hRvO#j
9 .��p8��c��¶Q�ڋ��=�N�Z計Z\�����u����۴o=��⿼����Ψo�@���$�[�C�2Lj�;����n�}��?������F�HJ� e^6�b���t�ڪ���ט�gu��]܍�<�o���4N��������~˕w���/9}�P��!��i37�W"�|�V|?�[�`��k���?��.�_2�V�կ)�o4�Э��Bp�{�p�B��-\��03�?�I
y�^��S$��n~�n6Vo�P��ֱ�B�9�i:�����N�,.#�0�����w�ڄOt�7��2)4��g\�'���BnK��i���B��~=����̽��"�Z��4�4荖���H�VCR���O�I�xH�Ӎ��z���ś�8����͛VM��@��x�qu��d�ۄ 5����2k�X\�������C�ڋ�yՓW(��Ǐ�";LTI,��㉣�N��s���@5?�ivo�%c��j$�w�;ժ�eY/E!6mN9���5���M_j?
��������|N1CP��h�5tL ��U���Q�ɽ"Yx��6�n|���a�y�&?�ޫWo[��O#��s�(��@�(t^����RT�x-e{��WZv��gc9dw��!�+^8�[CU����o��b}@^�P$�Գ(���%C� �!#��eBP���*�>,�=�̶�{1�ȯ��׶��qj[0�p�G[-bC4�x�8Y$�>Uot�-��RG���_^Ёp�D��=n��L�I̧ZĹ�*q��	�.~�A�D3����!e�LmX⚊L*"󌃕�.kyU���u�+�]U�Ǖ����x�V"A��8�q,b���C��������eW�%1�[;�`�ς�O���{އ��,=2ծ�ح:k�| ��4�=���ov���*��9������H�/Y�i���)���G��Ƶ�d��L #=P�5Ί���S�p�� ��q/��&鉯���ff�t�W6p�A����nF�qn�s�jJc�����'��	P>�T�a�M�\�l�i���+M_e]T4΄[.S@�u]�O�,hd2[|N��n0�Y͸�-���kB�L�)�Ǹ���?m�h��f�Wަ�,�����Ò����rVoi��#[y��xk�`��j����$���%�%�#������� ]A����g|�BO�O��jgS�ț����4;�wNA��a�n@�T<�O�!>#-�J�SpBd�2h�qM �H��
̎�Ͽ��O���!�o�<��e�C��&�n8h��;�hN90P�Ux�;ƣ�2�x������������ư�8ƅ���Y���O(P�˝����</}!ۊU��A�y�D�@��ŲD��)So@GS��\a1��Vĩp��l�`'�� c|���+*�<*�G�N�{̺<�1*��S櫂�/�ᙘ�ʉKƺ���+�D�N�� 7�+T;hլ�����`��:B�N��,�v �`m�����8��4�(���rխf�0&T~�+K�e>�p73-y�x����#�{͐�b�{3Yo�a��@#vn���"\�L�?Ų�֛��r��慼�[ju!Po��g~�"���"�8��SA�D�G�*5�ĦQ�Põy��&5���r��mX4�<ɢ
�*��WUbTc诶Q@*�h�UvB��'��zK~�]���^��$���'�# 8����BI�v_vL�t��.y4���c�zT���Wu���Ǌ��Â�������9V!>I7fHD�*��]S�^��1-���:�o�
�/]��4�Y��ة��>���~�2O�D�~��lL��,�(q�|bDvg,�B�3�*�q�y��=�op�i}Ǿc���4���|u>���)�|+��} p���������[����*�p.�X}=���)	n�{]�x���B6�%�M_�z!�����!�͸�O��4)���_]�����-�cǓϾ�8�`����ۈoXԤ�Lm
��F�p�츞^��-7x�c_o�Μ����u���Nh�����æ��i^8߁e(^O�"�������6�!!�i$�V*))��="��# H+R%�H�"RVO� ^Ϲ�𢡄5ҡoJ�l�����'��ce	���\�yH^��6�������TӶ�Xs���5�E4R����Y*:���jh��ؖ���!<_��B��d7�}��/C!Ǻ�Ŋ������������1i<����e����GCd���)O����8����j4�3���e;��1T�ya��l���ZTnLQ���<�Q�;��uc����|�).A��}�Z���2ȯ����}8or6�u��$]���
�w��	�W^� �`��z��Ӻ*�^ıe���� ��^�oĘ��)�?P�b�C4��{)N��R`,��}���n�G��~]�~B-A�ϕZ�\���X�62v�5�1���j�H�{_��{v��᨟��mQ/Ň��>ނ��p^=<�zșӶ3���а� �GX���rR��c����	= �P߈xF���8e�I��^m�C�v,؛��:��w���*L_82�ߏ�qw�G[ЎZ�{�!x�,"�A��������(�VGܳ�J�$�'�k����<�RO�[�9��z�p�3��WU��B�>0�*�ϴ����#�af��*z�֜���)_�+Ř\Wi�����dB��t���0�T�)i�_��A�\��bG��u���2�J7,�R=;{�f	0P��@�����|�v�?��m{ 6m�m�d��ۚ�T�H=��a��4�	Ũ�n�����܇��=A�A�wR�2J��:/���:a��n���%g.p_M|M��vy�������������dEy���Q��m��7�AWoe4o k��3�1����g�%�I,K�3��)��S���B�H�|��(�:��P�C���I������.f�k2o��{�f���W��4A�+�f"��bMփ�ל���Z�l?����F�g�}>� �xX�UL�Y>�A�'���e���9R�����&6JV@�]�%~���'�����'��RϮ�2��R�3( ��s@i�p,���aK6g���-�Ժ��I�?U��%�pVFe���b:�#]��*�ķ��bGcq ��7��GLjRް\�g ,�Cڰ��X�6�8�۩	%$�J��.2�7��#ي�����GfŬRZGd�pT��y�����b>��ʼ��wf���TA
��t�Yd���O}�(6��� �Vc��ӎ�Af���r�۶c��f�m\�KN�h�2�R\��Z�;O�(]��ub�Ԏ'����j�~�~!X`7� ���~W/*w��s�d_���A�<�-y�{������V��}l��?�5��X8��g<�[[���.>��m����'+�Ev6L������?��u�ϥ�1�;!���Q���;"P F��2-=D��b��AF�c�^G��Ż�F?��0�\5��Ȧ�'���T�w{�J�=*�8�C�>�����#�&miŚ
#|��v	��q��6
PW!�p�����EF�x=\ʲ_ ��@(������'ǲ�u`ܬ���y�����7�Z-��D�����%o�i||�<���?,}Ks�-!�+/"�F�anW�qa>0������n8�d&�_�Oswp[3�N�g��;v~��{��Řfo�=��:�*�x�"m�̷<�����򚠙� @􎤣I�~qPF�ȭ����5)Y�`ng�׳�p�S��Dۥv}��^$�����0Q�7�-��ɇ�U�X�Wƺ֔�7�*���0٥!#V�tX��
�ԏ���&��jř������G5=���Y�������#۾��M���S��
���&l����6>6�y�'<��T�_�J`E�Pc�F0)B�tbxYx�:E�%���Xڃ��Y�R�=4P�BN�-��&�1镂�#Ķ�¸����"�������j���7/���U�C.�H�v6�J�տ��^�z�����z��2��u��޲*�G���������[BA�6�7�����g��c�p���Y1�	X��-5]�ˍ�I�0߯(lJ���nr��H��(�'��|.��i�bk�^��'I�zo�>�R�ןWw��mv �E�Pi��{l���܂��0cV�����[�Ҭ�G�7��jp�g�j��^�C;&�,�(q��ñ))�^��a�lD�gH�z���#��B?b�\�����
\��|��eB�>�]��En��}��i�_y�9��SѶ7(qa/Q�zp��v�,�}�+�%#)��z���"j/}�!�&��q>iRC������k9�v�F5�u0�D� ��iBDg8���T�Q����5�%��^�3�QZ�rZg�����_�<:
ͭb/y��e�d�e������������_O����&�)y�s�%(o�a>+�o�C��!���ۏ3����7P$z;&|����t<D�F��n�.�~I/�'��������z����:t㻺�����$D�`ada2���2�4s��Ό�=W&���V�;E�Yϼq�ߪ�quѢE�����+��A�*�q�<�.���;����Y�e�a�\��G&�?Nb������&�
[��A`���lβ�L��+d�KH���A��d�(�#���h�P+\j���p�J��	5��iW�#��Ws�	(��m�J����'t�ΛM]����0͏�֙]��R��̰}��i�Y�
Y�ҡ�9�v��"��z! 4���f[�LX7�(��U�t��悪���ڹ)t2}�����ť �F2/�u�oM�6^΃k�"y/����&εZ+6�?�8�el�~�x�utQb8����A���J~Y�?�l�z♂����i�^��=��9�,\f�(��ȿɎ~I0�{u6I˶j��l�ב�쿲���.��t
��5N��á>}��z���B�o��N����M9fKMn�7�5�����>3��-��׭	9!�wg!4Ӟ��<ν�O��G�7^1ȳy^�L�U�����U�}xOկKh�π����@HY.ߥ�:W� �	��R�����Y�?���U��eƄ���6��*	�������t�}�TT�2�1_ZST��fWO�0�2Ҭn�d��7JRNY ���{|���枵3����p�ZQ�Ą����>��z�A���J�5���!�Y_�^N�kht�He�G�m�v@���*u�N����/�K �F�� �+>o�Zsk*�F��)�W~�Y
�� ӝi��;ƣ+�.S`���&�}�[�!��Ϧ�t���|q@ĝ��|]b�?Z�npi���l>Z�N�+�]�1�z��ܣ��3]ɜ�D��a$�c��uz`������!�czI�#��|,�1�#(@"�gتv�)[�a3;�U����t�#Ꮇ��)���ϲ)x�}ܳ�yx��]�|��`7�H�n��S�^@=LGV��رkR�Q�i�s�u�A� �K�"C�ע�mۗ��Y=�G�[S;8�&�t/�q�����p�3�?Jl��Q����&��o�RBҫ3N��I���I�Tá����C�3O���|&%�u�xfpG~�^Q�韸�ᠹɩ ��n9�����''1��p��1E2P���C���R��ɯ��=��8<�<ƨ��]�x�EX�%:����Z�$�����^�k3�C��x(�s�i��N%�	[�e;F�4Tb�b�g=���0��W�K�ɝ�(�X��=*�^G�F�>#0�1��m��|���u�'��5��	��v��O[{��+���%f�zImee`t��_�X�h3t�߹e8���h������4*X���d�vq��Z�Ԥ�P*vj*�G�:w����N.�WގpqQ����C/��B44���(��rf�G1x�.mcڒ[�?B�3�+?�r1�Ga��=�D����:`��af~K &`���Jx/v:���$b}����y��AQ�n��3]�@�<
+Q�$����hU��LI>
��ښ~0�ΚN4�H���lX\�ïP\�����*�����|���֖���,��|�}+�8�.�r�-�^�=dYEIc��ʕ��	����T7g������]�o5/��,PᏩ�ۆ���}t�H���u���uT�5ۥ���@�@���7�U��tr���` ��B�O��Jf�}-��� ����H	( �ح���#6��.jP}I@L�~~�犝�����ݷq��)�-w�I1���Œ�:�؟��ҕ��F�牎�0�Rg�����d�����@����i���0���s�0�J�!�91#�}`�+��D�\(c+"��}GD�8�nh�A����f�2?�}���)�h�]��8}�g�@�El{s�b�kL@i�ҒU�V�4�����&�O���[�rBR͒��VO#}pN/p����"+H�A���猕� ɡ��F�n���&�<M�2��,6T��K��R�?�Nt�	ѣ��t��cFJ���ޥx�u)�zЅEL���|������9~����NJ��/���8 �R���<ְ��|/T��UzP�fIѝτ(|~����'p�&���~=����R�vK���Zrf�ڭI�����%=7�&!*�'	��W�F����:2'�(K��6A^�!F
���O����;���Wؘ����u�0�c%VJ_?���Y��e[��]�	���tLD�HJ�j�"A3�jMH��Xe���C�qW5S��-!-�.\�\������ I�cJ˗.��%�s&���~S��ɉ���l_���9��QhaȔ��b⤄|L���>k�s4��_�^�ƒ�Υ��`^^�F
I�g��,B�2֑�	�]DƗ����+賗X0�mC4y�f;�/�V,U�2k���3o緳2#6	e)�����!2, z+� ö��:�`cG����?񒳇@y��v�(� z.��D��ˌ��Ŕ%�����R���G�0�'T��۟q�v��~u`� ����I�X,]�&'z�Cd�2[�r����:����Awn�p0`�� �=Wn�K���$z�h�{4:\�f�C����{2B��~�Ь��j(�l�;#�U�\���D�h��>�=|�"�[���s,���X�U#�83��M�Dm3��R�,�-keB���uo�KjW��:�UT ��5�����-	��Փ�F��Օs�q�{1D���6ǩ��NUxO�Y�Rr�̿�� ��v��RZ_�fz�8�Ƕ��mzcD%m���o���H@��#�g����ޜ� ��W���b�C��I�q ���v%k/����W�6��tǘ�i���HY���K8@&�G�����C�A\r��0%��\��$�V��U��c��:ƃk��3dR��<h��4��U�d�F��&Y�^�(�t�k4���~�s��Τ�����6�v�.I`�]�C��&z@�6H��]��,�PM��#$�ۦ3o��nE���Cf�P?.݃�% J��S��g1���Ú��{��'��\�ea�%��Ѻ�T���|�������}\qO璑 �ҭ��bʩ��0O�ZB���I�nl�:y��x95�=�Q�s�@��U΄���X��1 K�����d��Tm�()�ǚ
�^�(�Bg��ف�����"�(��H�M��JMf{Pe�u�-��k��0J?ԡ��;Y��_Ƕ���d���$��(����^�R���7+�q-8w��W���\^��\M���`@P*�hݭ��?|�
r��^��2�۵j�¯��7HJ4��xj!�l��m��4}�PǊ%���� �|d9��I���W8�κf��j뚧���G�����Q}�ֈ��
�w�Z���%Yv����w 7���&"�ӗjg�l=vЊ����Oiڪ�ΕkF���i]��qB='�M\?���Q�bU�Nv�+q���#82�N�KZ� ��]���~奙b�-��<q.,t�<�>ב��W�M�
�5H��E��ޅ�Ye�H��qM3*�>OG6������!�,�:�ow�&�v<l�����!S\�cEv4�R��ҠZ|��e��#;�,:"�2[�Z��u�_K`� άU��G�'��8�g��ݭ�"a�[	ʐ��'oj+�M8ddW�Bְ��pזK{Yp��#���'�[�yg'�a����M���h�ИJ�;�����#�
�_��~;���kD[��U��B�-!@c��>P���K��jyJ�fh�|����*�ֶW:��/_EGt���?9�ƞ��L�#
�������	��8w2e�T�\}-fET]�x�[�h�x��l'�b\�L2����0�����ʞ�1R�P�h�T�H�I�����x���)�@�1���	�sՒj��5-I��
���@!�Ȅk��xG
�\��_�c^B�����՝c�e�@z�9M�|�ͮ���%��j��$b�(�6%�ݱ�t���*������d�|�&�����^xLҞݷ�9���,�]z�jZ@�ᠵ[Jf闈MPx��"}uo<7��7L���"�$ ���zCL����=\��b�	���H�y_��a��R:�zc�P�XBl�;���HЕC2�eY�!
�\i�)�#!����I�O'"7��H��g�@,sz���h;=Zl7�����>�?��][[v��5��d-�{T��24��ᣲV�&��%w��3�+' !��?��ۇ!
�_t���oT�3��hY�90�B�\ҵmD���G�m6�Ǒ*LQ�^&����{c�� v;�w	X:q��T��*M {����ҟ}�*�
�8tm)1Q���$���o)����n_<a{�at�« ����2��=����qW�Ӈ�>0k�43秌�Q1���
���{�[��bI^8W�v��?OP�HbT27Q�ٞ�99v����.IL63,���N�<�71��-��2NE��0];Jc�\��3����}5�ݞy��J�Q��_�ll�9m�|�b�м��C��g�@���J� ^*��+uah�ǁBy��d�aoSCn&�*2����W�d;�19'���p�D�ƣ��,bC�J��-�@(UǠ#�ZCpt�~1���O��Շa��Ɏ�@h�6֭�<=� �L���դ��df��Q���F�^��ۦj.=�ג�/����o��=�WN╋�|���ΌK�A I�Z��^�ds�����Mx"㪑x�L��&i�G��K��pͻK�R��|7U�iQcQ�v���f9�b@�n�|a��AjS�р3��[7�-X�cw��p�}y����$�����M�َ���5��T�z�B4E�*	�}�9���#i���Z�AW�~g�L��ѭ/%'���n����G����R@���l�f7�q���2�Ǌ�f�q�:u<Rս��9u�c��m�s�IU��9��ꭸ������FpT�8S�C�*u�z�e��qHoƴ��㲰ћu��Z�װ?��S��D�s�-PQ��+�����s۲�$8�?�ȵ�[��~�@�� �����vٚ�����X!Xy�ȫ���%�D�򓨁i�3�r{�N+��~���ֱP��
���!�Bۗl�'�zLM��e�D��2x�,�<�����'z�Wg/'�Ƣ�t��5���.����o�;H�@�pbLpy��km���Ez�6�d>��ѣr��.��ңt�r��΢��w�ң#�'���f��]'tu�?I��@���v�wȍ��.�aX7�D9y8��D����"��x�����vO��DV�/��X;2�.��4���$�{�R�y >�%ǂR�Ps3,�R-�A�n� ��%~L�E�H�̑\>���>(���k���O����Z�|g���R������MDI�Y��'���	���Gی;�2�|Ǐ��۶U��:��� �:sR\O��NbO]ٛǘ�s�)R�*���룇�Q�+�{̴��K�BA�+r�تh����m��i�k3P�h�2� �x 4F��P���$��H-�$���sփYm<1���k�c@�6�Ǆ�8F��N�L�N˙+p�1w��b�wF47�|�jUX*i�.K1 >���߭
pB*�AQE>B���HY������-�#�G���꟟���m��h8Jcsym�� S�K7D�o��)Uo>��L^�W��gȪ��.�	�x�~8�n�`uPQ���7�5��h����e�ܷ~�0H��#c�QDk����F�I�N[��6�\�T��Iw]���ƨѷ��T��1��B����;r�Q��M��zĴ!�3��s��E���P��r�(�h�E�&�B⺧��[�o���2̊�V�-����� �_+�i5�P8��Ӛ����`QU^���]���:ƊK�G�zr��MwW˵�>W�N����}�lm�j+��`ۚ��
�������Q�'i��a��ϴ@���W�¿B�$���F#�������'� #г#A?jg��ul�ײ������⹭+rl�1�c<��� N�=aSVдjS)}I_JA�<ߦ2DI�$���ل�-��)�ô��C��~u�Ѕ�#�s�(6�ir*�%D|�iDl:��\��:���ڙu�0㟊�՗@mq�¨CI{2�:�ɷ��<����u���7������=H�4*��/��U �Ns�,� ���z�vl�'�'@��EtPI?:�iܬ�7���ܶ��m,RM��`�£��~����C�q��`O�D�k���V�_0?�7�,?ڪC*���Imf7T<P�Ԫ���6`Ak�g2���;|� K����5�~�"w�(��qh5��_��H�qO��e�Z�J�D����7�8̌�.�*?G-U+ʿT�͹!��&�l�~n�:��������t
xr~��o �]^oD���d�"���۱d2ü8-Hi${�̆��yzn�ma������x>�I��.�fޒ�[E��_�u��]h���E����PY�v����~M�u��	iOhOH2��$�����C�U�j���$D��I��/��9.�ҏ2�u�X���Z#:��_>��l��U3�S��]ɤ1��s�6B-��U������9��!n�.�*�|�)�h�I��@&�5����D\�h��}|�7'lt�H��'�����'Gp��der+����4O��g:�`���E�\������C*��`��x,�`�lq�1�_4A8�[>������`���Ո��f�Y�����������j<h����ܘ�ScI�Iw YHH�K+�F� �‥\��9����r��p=Y��T�w�U���A�˝�
Ɂ(��*o�V��ʯ�1VRC�b̔uG����A����-A׾V��(�P���d�Ó�k5@��T�0r� SS�U:�Tp�A��~B}���G|�^-~2*;�CV�#]���ʆ�o�qΟ���㗏W�FA�љS�r?����0/�;?�C���i[>H]2z{��W}$�:�O�9���s�/f���9�.�Xy��8��K'L�������3����R����p���C�O"���&o���̄6VΒ$;j���`$uJ�>�1�~���!�3ri~�ES��Dn@*4�X>���������o��[j��5G�ߓ����/�1�9DH����\�8`&�\� �E��]�M��Y28�Ywd�S�n����ypOz�%wh�ڋ܋g��P���c��Tr����g��ǖ$�����/\Ѫcm��%8�-`.;{������Ĝ�8������=?�6�.+�c4�y���N���K�_��_bj�&��`�l6m7X��QL��c�Z�~$yW����!��=|�Z�W�;�X*�U�y�����L�\��2�&���	��##���')e��"It�@�ؖ��a��ÅZ��5�I��v7S�:s��أak�K�qҧxA��`��"���r��5䌣�2A��#���r�2�M��w"l�j_p[
�l��w#cN�l�q" �ǩ��k�9e�`k4<� #�@�y� ዆�{8UD���$�˃��Z�5��*���R�B&_J)R�C�n�٬ۤZ�9ҿ�e���@\+��8=�$d�o�ZI5�my�C"�ȡF��%���C1��%d��'�(%:B��x���ϱ�K(/($ټ@���Za���?�Ye��,݇L�RΠY�^}g��O��?+]�c��OB2�Z�D3O�p��	D�M��Sm0H��E��O&<S��� #�3�D�3����[������ʡ"ֽ�����^�'&�|�/>����F��$l��Y�-�P�>��&ay�$w���v�ɹ����h��M|�$��S������wo�N��<��Q�.ϰ��]�Hd��0��Z!�<���4�	�$j鯪�75������q���f�V��xO���ӊ[lR����8?���z1�r��E����$�|�x�{
}�8:��U�=�,G�˅n��%�p��P�W���/:�@�Ն���2x��l���$`�."l�f��fN����"�$�(>���f�ް}}�̻�]�[�u�\��j�!r�2>"5ٓ��CY�N��L�j��VM�l'm�ܭ\�hAΓ L��T�ⵆ��dO��e��e+�E����Z��vG^�P��i����m�� `��4���ҘI��7@�=���ù�9K��3���2�BEJ�+-/����3�~_�`�a
��p��ֿ�
H��AtY�js@���;'u�~	���]{�574_pDXʣ�sG�z`�S_S �;����Y�,/��\;ǟ�H��u�h�(��M@���(<u�m�Sä++ƥ�a����6 6?r���g):���p��G���|���E���͏l�LJ�>��8�����9w7�:�+�X
�A��>z���㮉�Y:h%$�}PY
E~���v����ϖ�������î'HW�`� ���Ep�� x?2�&ۃ�����p�$��o���;�c ;ި�#\d9�T܊s����ӑ�Fzڋ��4�~��0;�_Cd���
zWO�y�(�ڄhF.+4�hW����<=��a ,|��P��=R��x�l�_��~T}��Y���e����׏��Gpn�,~?��#�Ϲ�6�HIT`���}�T�Pt�;�
W���De;R�1��N�~c����i:ta Y���W��X���dc�R���=�[�jf_�M&�Hr����V��jb9�rl��~�?���}}�%S�:�B��4��{+�V T�k�����t�BB~�2�%�����1�q~8^ބ���JL�/c����0a���t��ȬB�I6�<[�4s�M]�pha��59����̬^l6��9���\fk���_��}��;A'%�d#`�e�'61��W��}c �g���\�6�����?��4`��¬���wg݀ҿm�
w�[W3�ɰx�:��;���%�<$�Z��Qk�P0��'�G1�W�K�ѕ3���݈�pe@�$��nR,$�yw�Â�Y�K���w�͋�ABn>�͎��ì��GR��C_E�8�y"ѓ�,�	�ҏ���"��͙��� ��H�A��z�j��ư�i����Nސ`1I̊ �7O��U\��s4�=�ކ�������%7���>Kg����3[�=�ĥj�)�~���ޓ��5�}o�KeŤP���N��_E�g��I���<�&���J�Y�}fe�ポ{��!J���'�W<���Oؼ�I�>����o7Mz
����K�r���U��
�F/�"�ӓ�|�C�v�1��3��l��O-SGP|g{`1��8Sj�Յ^lٯNɇ�z?:j>h��vފAˢ���XHG� �F�Lv����I�c��'�.��ɾ����С�^�SjmP�j�O�����qZĘ��t��X||�(f����7����:+u�7�2���|�V'�R�3��$}v�BV/�w֥��rRt'z�r=�����"�`{?V�ZC
b�Z��ؿ�"w�Ē��"ùS
�oj�zf��W�}	�U�v���܀C_��h�6�H��3�����������5&>�V��ύT�OWȴ5�,����t��x5�ބ�̠W�ŴF���YL�ѧ�yD��� ]مv��±� e��?���������%њ��J��2<��G�"��^�ŪHl��]8��X��gsX-���M|�x�l�2�(q����P����gi[[6l�5�*/f�G^�G掭O38�� X�����
cz�ֺ�ɾ�������-$4�=#˳`�!H�����}��Y7n�����Jcq�yz�0���1h�o>Q�O^VѡI$�D%~�\d������[��6�p����,ޯ:�{ �-?��x�"��摮����5��@�Nh��^w���DW�Џyb="e���.iM0e�l���`�
�J'�g�ݘ��d�% E��n�QL0��MRSx���� �����L�f�,��G8�wQ�o"MwE1�pd����z*�,���O��4~`Zg�3�?>T� z��w�ᖀ��\�e�BE�.LH)|7xk��b#��EG�-4�d?��".c��6���=4Q]E�sN��~�E2��\��D>� ,�+�Kpt�v	`�ЕI�b�%,��<��[���`�Ԧ~�j����0��˄8��Ҍ���}���|�2#��b��$���mqת��K;�.�Զ�+����`��
��-�P섉)����-���Z��(�:����y_6�Ւ������+�ƴ��n�s��U���5!��WU���]����ڲVu�������KHoZƠG�l@^����M{���Pvc	սR�m�9��\��A��j	4�t0��m���r��=��X��vr؊�����Eo�m����Kdm�j�=��U����"��4i)�< �`ukZ�F&oI �b�O��З�-`��i	���
(��[�$cQ}�q�4�So>�V�C�>���p�7_z�J�,E_6����t����)WZ�Bk�m0J���]S�ڶ벝��{U-Ӏ�bKk�������Iȏ�iA$�)m��]�ފ�0b���ɤ}0e0"b��[�&s�x���6;_b�����I���XA��a��.�_�Vn�a�|�8,��
~+H�}�Bڤ�?�v�$r�>zu�M&��"8m�g�<�WV���-��_/�]M?�|ԞJ/g@b�F�G�7���l��o�Q�Cb��#CX��Ǳ
�.'���W"Qu��4�?�r�i��|�6�P��[�C�u������F��^�#T�]��[a8�	�E�F�k9�����HT>G~���"GY���*k�v�Y�ֹ �v��(�9Q�����I7E��ڟ�Z�����M1s*�}˝�E�ss��uU�q	)eV�MQA'��L|�D��s�ai}�;f2�������	<�����h�qMƜN�+ܝ`.�*�f�s$�a%9�<׼����yp�6�20���џ�D�x�t��Lz;�CQ<��݁UZ#vD�-�h�y�}no� $��|���<���*��(��@l���2Y/��B9נB��e"2�@��.���������bLd��)����q��J�Dx�q cH���-w0ɣ�nY��)�y��ψ�]�{1��T�,/}Ȓ4�??D/)yh䳛�[q������W�ƨ��-��mŷB�ԏs�]�#�
�c�m<�o�����Gz���h�+�S��ح���p��vpPn(���묓���N\|A�f�ٴ#�.kLC��5�$	m�?�a�����Д:��XF�)�G�l��	$SȔr�Ԓ����'a^r�1*?Y�2��K�r��=B�7�(eR�O��-{���Z��<U(e�c�b��˝0��[�}���(Dh�r�R�v�?o�V�[#���T��K"��H�q^R�~0��6�:��0a*�ٗ����v��jyocE�)4�؍p>p�5�YY(��V�8��p��[m:FxN:�*�B�G��|�@�����G�!4�oDT�C�?���Ѣ�D$Ug4�능l\,�@8A�%P�!�͢�s��3�'2���A����f�������*dQ��uB��T��L)���n��6�@L��Sv���h?w�~-m�Y354�<�lb�)x��|̭o�}�Q.r,��U:�9���IQW<�8W��*GMr��h��G��'��ٓy9�����X�	�(���s�
Wa{W?к6_�:�Jn�*�=q�W-׿\B�&/�)Puz��m0�B�@��j�w�r��X�F_�D���A�3��H}Z�0l�T�������{�B2-[v�P�Ն� '�H�D
������ԗ�O�����j.�&��ĥ�eH,(]�\>��_H��y%AsU�"텃D_��ڇ�1�މilS&�6�rߙY�����zDs���^b .�W#������Nh�_Pi��ʟΦY
ā_9ϩ�Y���V�0/[���F���^�/r��r�r΍^���-�03h*� 	)�w�=(�z�W�� ���{�f���|�<��vM3��7Cq��nmL]���AL��G���1W��A��'���N�Ur����
��sșpe�R�y���CD�y]�J��cna�����JfB�6%�n(/d��m<��B�`��}�{I��*�a��|��k"� ��!e���N����!~B`ס�tM�����{�\/�b��Jk�fnL ��DP�ˆP��9����5������$�RQd���8����l�$���of�=����t�/+���"�l	�;�RW�l�^�i�lr�r�e��TJ-Z�_�
�h⊳u%���$���TV�y/QO4��^C3���~����g�՗v#W�Bk?�@���Dp���(��N�JC�o�I&�Xv�o
�.�ȕ��)��G���y�#����=�4P{�B>�ʮ����4а��<,v��|U���u�%b�m�_&ʃ}Ȕs.���҆& 戄;d��n�x�<S�Km,�C3�t4�gˆ77�����B��In���	 �q�U�8ĝv�P{{	e3����D�~���aQȺ3G�� �D po�s+*b��8#��tr��<�MW����)��ܺǐ�b��i��mB��_�	kzv"�?���u˼��փ5��,Q�l�s���4k�j�Lu#�d��4{��	���� N�3c�ˬ������{s��u[��׎�����Of�X�Q�!��O/�ʈ1v\7���o�.�c���!J���%T�]L��p�Y��.��Xȟ���d*���U1��;�^u������A�Z�L�En}7`�2I_9��|.���k_Z��"z���43��ǖ0I�e���m��1�O��������Dc?YQ2A
ye�l�%��� .94|���aP�u�vHb��*(��w����*a3=W����$�B�e��Y2�1z�Z��y#>���N�n�W�F�IVVD��	4O�%'�!�����o��}�&瑽꠶�Y<�8r]+�mꅪ�Z"Yx1�ٱ�%2�>��������]���k"�6�lM wtnT*XK�nՋ��R3���o�F����K�/}	C}ѤX-l��h�idB1>��"PU�%����9���������6u��쾯�����Z� u�6�JTX��^��e)ղ;�1�?�5�*;d�\��#3�-	ګr���nW�3(��r	�t^"�1��dEx��b���Še�5# ��LN�O�vܵ���7���dw��h	PS���o�2��i���K�Ǖ����}B5:1؂�.O�aw��^����8�:��$e�׀̎�G�}���	��L)[c9؀퇁��L54Y��ىl�
��伓�tq�³��8D�@�����J�V-D���"��I���7���(Û���_ۭ%�b3za�6�fq%�������	E(t�xʪ��/+���fq�m׮�r�޴�C���^���0������ȃ�a`��3Qq,�tDA�ǖ3�@��X>˯���M���y鿷(_���>�uQυ�qz���j◲,�|RA�*;lZQ��UT���)6�L���ڽ|���5k�}�j�{숫W��I'(�����<�~��&����ѣ_��m�8[�k+���+lwT�C���,�M�K15���`D@l<�s�"�ݝ_��u;����p�5�����#$�]lu
v]7���>��@� �CL]�*�Y��,�|��˴?�$W�F���hϣ�db�I��D���ܤ���lA�ǟ �=�_k�,fo�(m��Pg���.6 O&���M�J(D5v�M9]��[��".Ʒ4'�eЛ�x8`��F�=����%55�6�d�=����j��N�˴��:tC�k�8I&�>Z���Y�L���\�x>-V��7�L	�('�osi�-��]j�q�B�f����[�K_�H�e�a���}
�&i�~�M���6�$r��4SA���'�L7�tdD2�Ϙ���KE�����ؙD��]���+��*gz��;��z�7kvr� {�ve��o�{*X��
�s���}脡�Y�x��-���!G��WBk��|���{���۫~�M��p���r��y�j���e�d"�-��ؾm���J��=�*�����>��AܱKV�zn\�@͏��U����C�����9r�0 �s������)��5������f�\/s���5����A˱c���w�s�J�pB!;֓{5�E�G��~ ��U��ؑ���`]�|���sYHz�'Ss���UF������a����/Ba��ζ���WEbD&qBHSU��S��P�1�K?[WX�]�^ ��b�6��1�jc2��|Z>�xo�+�䢌Ĵ�[(��X/��T��Է����,��y�Έ����43jxx��*׃�D)P��r�A�d�t�ᱰWy�pt^-O�|&w7�Lצ �]ئ$�R�Fw�@�c�*7��eYI(��چ��������)`A������ r퍾Kna�"O{��+B������+�i�mH�1L��͓��FX=Т�q�����Z�P�0��M�e��׶W#7lO�������D�ݯ��8��nJ���:�۷j�9��C3�n#�D�OL�ۑs��Р��N���>�(i��&Ɏ�\<���T�fzV6MQ�cR�%�u�� �&*.��SW��-�;�I^ึ�&���u&�1�B�i)�n��mB�$����YY-	(�������\��'ӲB��.fkn��/����V�tXo������B��pزtٽA
=�_xØcM����J�Q���Q�N���~{K��=�{��
F����������H:	y;�e�g�K�V���u�1��KR����)��q'|k�Ut5�7N_� ��_C|�\��κ�O�wT�V�d��e�*7��-VK�3��'�ѱ;X]���cۃ|js�+;\��N.�{��q���F-����D��S(�mD�5T�������u>N;�К<1MJ��o!�Q�'� �Ev�d�m������D]D,Y?N���a5/}O�R�,�4�k����j����s2z��Rc���I�R;V��u7^��3[���Uz��� �Zԗ��ۄ�>��>{&���<ڈA��'Zw���<���4��&�w�5IusE��ㄘ���݀�^��0�[^�s���\�x�����^����%��wi���)"��*)�j��� **�7��
�P�+��1��4Y���K��Xt��t� $�(���`x*��E���qUiq�H��=�g����+��o�f����~S,u����)��3;fcU�Μks��QлB�W��X��{����$�KyB��=lP��)\����ڈI�$�1{�
�����:�+�ւ�'=2S���"�q9������E6#��#���1��ʯ���ڳ��"qڍr<��n_ю��i�����Nr}�{=|YV�󴘙�&5��>d"�p��?i�t	|*�I2�	*��j�w?2v;�7���E��6$�]�]�݃�B>��f���Ϗq��8����'�<�պ(�!Ԏ2P`�������G?BC�q%oI�e$1�i����s��B�-�&ɢ��] d�eܴ�/��ޘ-����-)����/kSB�\���~�8w�����{��*��(�$j�$��}^��eBT��^�(��̰C6���H},vM�/{G��b9�|o�����8s����,;�3m��h_gSv�jm��jX3��:�������+�B;�Y�p�)����.f���բ㽄qwb9���sR JCj���c�����%n�_�N�F�
�Iu�t^?���)�je�\����L��=���΍[��D>�Q���VM���M�1��Xp�e�ˌ�@p����B=2�l=RO���3##1��E3`�˚b���ob�Ԝ����w���?�[XrŖ�|kh�_��ȟ�i�5$ vQ��ob���_�A���o.�i�kFLe��1i��SC9]qV��r;��7��H����rX�w䔖l�Ev�]Z$]���
\���x��)= ����$��0bD
icJ�u�}4��AYٓ����� ^C���d�e��Ū� �M\O�#��ٟK�m���B�Io��_ �Oq�,z݆c����F��F(�]�F7.�o���YM�Ǐ5�J�������W���;�u;t466���F�2�$���>�$� �T���L5h,�_\������2d�R0��4��y&"+�i"yn��/�Y��	�(�6�Q���?�ݿ��	�X�"u�e��hAq�+�j.���|�̝��3�'��tn+ȊrՒ�Fl�HvN�8}C����J
�JzKFX���1),� �H�Y%�ĊC�Ɣ���{i�a~���엕b���	��Jt�$2�����!Gb�S��)��7�"Mu6y2k��k5ztڐ�M��r�7�J!z*B��_�y�|���;�c��pi	���[ݍ���qx������U�#�+��:2�_ɨ�ck)�bh�F&����M&�1�3"���.����֋����$�~��M��@�L���1nB �RI��8���Ɨ�	wIž%��H�	R�"�I\S�xw�a����;o(�-a��(�Z�������#K!A۲��C�e*6��a	Fo��]U��մq��r�h����?�]qB�N�"�LQo��0��M�8jMn���^�|<��Dj{�E%0����D�{Y��ľ�#��׆����d�5C|�� }����u2�$��BDT7�id͹|�}B���b]5�z�~��sB������� HgW��#���B�����EcD����1���B�/��>�2�J��Q(��%��D$�0ٸ��L�1���ZU�Zd6k�|+�3�u���ʹo��?=��O������7�-��](��
'7]*�@d~�qF��C˚n(D�Wc�7UH��[�vNk��^�$k�С̛Cκ0Y8+�k��+����f=4�Ծ9��s u���ղ������_�yu�<���A�=�����p��*Ჸ2�Խx3d���;4*;���U��R�g�������2aiꦀ���r�7|-f\�w�)
�Cڹ�����2���9�^���͍]Y�N6�W�"��m���]c�$�/8սW����lk�U����¿1�<WV��,[�۫�ɥ��>&�H��Q�S�<ΗE�<$��؜���/@�\��J.��p��kc~�OQ�;��qRnצ�ʟ$�2����J���6;;v�H��-k��6��eO�PD����$N�WP�AQ���,G�W���P�z4��v	퀘l�W�y�ڇK�nM�ފ!���~	��y �1m<NM�R���� :��3.��0��f9��fZ.~��L�btXu�f��N:3}h�GV�4���`��,v���>=	���(X�?��Ƒ���2Lz;���׹;]��4���;+��yڀ�J8���>� a�@\Y{�/��m�F~�hMX�X�a[>��:v`Gjofe�a�������l���R&�\��%+w>҂+Y$�z�0Y-�?�S�7�.�^,���O�ޗ"LL+VA?��ے��D�Z�֍ ?��lt��i��J4��OqX�~h^8�|��4E3�:�e�B��j}°���$̑Ѹ�M�r~�$�g�f�h�@N�AKh[u�zötvy�!x��[�g�kK�ف�}�KCH�*�vZ\8��hK��7#���!��O0ٲ���)0������īgB#q����O�80��4��6��HW���w���B<d�bF�Nh�7'S���N�-#��T��TnM�����U��8��6%���8Sy�N��؟��j�&��;�����kĚ�
��G�m5�N4V,�X��FX���YI�ƪӀSr,މ��n�w�j����蘶O�I>�`���_�R}��&A�S�J���P����=�̠1}(���.�_]1qkL�U�
<_���Ϣ�n�n`ɾ���7�-ϞjF�����_�M�T͢���dI�B[!���*	#�[����yK�^5�e9W���1I-스�H�OX�� 蘍]��&e<n��v���C��*u�o0"�(ʿ }��F�ާ�B���mF8��_x��3���&�	�@�˵�(���n�I�����L��$�iMB�XIv��b?@��5�^g9�`�C]ㅊU~�WH�n�h~53,|/ڠO7jR�;_�&�Mp��9���E'fI!� �gY�{vX���)AR�o�'5_v"mY!��$6c�à���,�U���Q�,��9�{&��'ҷ�̱�G���Y�Ǟ����aS�:ӝ�}x����"6�_�_g(|�=�m�-9f0�!SQ²yyf.���B��)�����hn9�
e�,_�����}�y���fG��4�����[j����"[�T-�qM���i�y�>����Fo���_@^�>H;�����I�^�6�"��Xp��h���v�+���l�R�0Y�	Y}��Iŷ��35v�9�������	K�����9�0�����i_������P���g�Ż�o������孧�Aȿ��ۥ����
I7f����~�,6�)�t�TT Y��k&Oǈ��,�x�(����\�\�x ����ꐕU�%'�m��X�
(>0�2[�8nXSEp	����.�򨏹4�0v���Q�0n�u�(6B�s&!u��9��̕k�U=��G~��/d��p�[Y�kgTM�+ks����x�g<#e9�u��.�{9������ꋮ����l��<��?�yu����a��	�'7��Ϳ0G��K����E�9UR9��c�5�r/�\�a{�@+�mٟ���I�w#<�;��A䪰�'�����I�S�65i�R�Q������,�ٵ��\���ɖk����Y�^��Lq-UA���� ��#,�a3����+a?�� �J^H���s����ݸC�_q��cA"��)�M�J�73tB䥙��:`�8%綳�9��XA�/���YO"�+F�K��&�UL6J�Jzl�~�y2�v��8d+���*|ڹ�z��u���J[�_�#�!�7@����:��+.�v�90����m��Kq�������m�>���Q���},�e����[�c��%�B��e-��=�>*��x^5��9vZL�f�]>�)�> � ���?��P��]2��o���|h�̉	�����1�0sV��$��r���]B �,jk��*�f�M-���Fu����I��,�~����V��;�۳�YAĩ�J|;��Q5�n�DU�ծK�??�
� �\�N�l�a	i+hql�v{�{���-�A8�oΉ`�5�T\��*j�ܓ����1�����`O԰N	w�X��\�ܦ��1��^�<`/�2g���|�Z�=5�A	�`�	z� z����o@�ټչ�8_d�-a���偑�7~^���E�Sk�`9;�s�uX9�.iYa���~�X�|j!��hc����4���=�b��]%M��QGe��O�- g
�Dǹt���C�c�Ϥ�`�����ЌÏ�l����S<B�E��.����5��d��@�KO��P� Y���Se�����NpA:T?�㰻lj���܁�YKM��2��m3:��=^����*��cc	��&�]j9�m��{�/"�/:֟���˩�H_���?�T{, A��.��t��l�g�=&_ O��Z}Qb�/9 Ϸ��������8�҈S���e��7��$ ����aE������p:M��_��US�e|8[c�(i����#q$���]���K�q�Edq�Q�  &Ц�{����s��n��ܭ�Å�����L�ݢ�-��THσ#�>Z�^���B�)1�q�|�>&`b�������+Ӈ
��R��X�8��SV�â	)tl����?\�b}�����o>������k��+�� B��=t�����^/@r��2�PdR��uPcj�s2��ױ�+�aPk��վo����>�"��ca=��p��R��&ۦ%�QC�����kr��Z�1f�Z Y��������D��Fx�%+4`u3���LC��]8?f3���~ȧʿ�q�S:e�m�;u��a<R'H)J�2-}j�� bz�?�#.�0�v���-l����7*�#�R�i�ad@�=��.�/�&-Kr��5A&��-�D�n�SGtm�1�/����� ��Eob���7��!I����;2ax���h ��E����*3ʜ;����������ӷ� �!��ш����H;�`
g���Ϲ(b<�2o;�n�U�[����b<��4��څ����-{6�}7�a݌ȄP�:~�|��"N�����i�E�G��:����e�W�2�ͩ��mL�|��Nr�y|����߅�S�:�o�"��&�a(�oȂ�ia+�ی��# ��ֳ�/?.I�c���ރ�ƾ����m>�*�&�Y��r7K����n�� >s������������K�Nv�N;����>���=�
�i��?F�O���J�2��NĚ�a�e�m�����#UE�M���|�Wj�f�q��4���q��ۛΕ�![��YM��܄%�r̞���Fj@2 �.0M�w���=fn�T�}���Sz�{�z\/B�,{�f|���,8P���n	����$�+�{�%1T�4<O�D~Gy*�$�ʚ��7�2�I�]�jń���vG�}�:Vǋ��R#�pXCyQD.���Sq��2���!1:�C����{����*����ˎ�q���_;`m�ݻ?�h�h���+UTY�]U��_VT��9��:�}����� �'Ẉ�s�%y\�C����n���c\��[.�4�P�CEx�"!�h�4��歂�cX��>��{ F��wgy �'���vK`�CT8������4�˶�3����ec�y���^�ݥ�L��[ s��M���O�B��)�M����8�s�!��U�j��ʽ�NX�����$�+�b5�2~
7|����Ke�ߢ*��JM�鯨�|F �����6���m� �dӚK#�[��9�˼r=�	� ���f��6�gQ/��QT|�=T�ډ��R����ںʼFqSt�L�]���X*p�4��
:�nh5�&t�M��ҩ�8���/�m�\�ٟݎ#�:��h00��n��ݚ��J�`8���Y���6��3�ՙĤ>�fk��@G�j�>�%?b�@n�\����m�H|e�siku��dy������:��p����NNal{�1��~����PhJY;?���]���d~��8�N��yBϥ���T^tb��bBcn?tޙUU~ƂH�)������A��w�) �N���]<륯�
�JCS��7	���Q�YL���]���XI��[�	�qd���W���$�`��?B��A$��o<��[���@��D�����[jO�L�eU�Z.�<W�!~�:ˉVw���ޔսp�a��I6�jkH�4�|�<ֈAy�Լ��Evw�u�mN�� $����S#oP&FI$�.����ܧ�8 �g���i�T�v�Rr;J��Ѡ�R�Y��r-�-b��^���n$�ؽ�?m�(2]�@���N�v��~*ԉE���x��b�H����I,��dt�C��K�/~3��Q'$�j2g��t��_3�6��h�,ީ%d��4�l;=�X�\�
�2#���tXy�n�W�1wwېn�m�tSҝ�J�i4�R�j�V�>xM7܌�4|7%cp�ވU�bZ)���;F��c��jW�{h�v�EJ	TF@���V\S�����:֋Y���]^������O߲�j�<)J{H�FŞG�R�.�)Y{�ck~��;�y(�|V4;�y�g��ֵ·�}E����W��-��a�f�����;)Z&S��(W��}&�?`~��P4�E��"΃ܣu��,t���2v%�c�t�k}��<r&���˿��s(;�Mx�p��@FRX.iz1U�{X��<R�5V�-�7@�P��C��i���$R!���Y�Fi�l�j�CHѩ-:.�<�΃�}�z�d���"(6SJԦ���p���1�{��k"	x������#Xl�����+�Cd��:>�@N��wz�C���Ցk|�1r�����?���ǭ��/Ǉ�9+:t�ؒ�4Tz�2(;o��)��c�-�p�S�qL�]��='�{�v:�'�ﮌ{2`0⿀a��eޭ`3��Q�{�a�����m���6T\mpZ\79bd��3wd���(��K�͛"�U]\zPX�7�|�Ꭲ���m@�q��o/�qX��RyK�&wJ���aV �ĸ%�� ���mC�0]\�� ��3O��hv��_+�Le�(K	��I'J�f-�✙N� vY&��j@o)�/(<�����D֩!����ߔ˕[�-���lc	�`��$����� ���_Ý��,�����1�����(R���A�R��zs��G��l��g�_�%�f���N0F-x�$�^W7�Ͳ�7��d[ZQ�0�ܟ�"�,�v�Nl��j��I���k((�z��Ap�=¼�]�1�C���zVԨܲ�rQ|r���J��lހ.<�&	�r�&l�+v,b���a��v��5�}���SEx��G���	@��oP '�r��cM��D,ˋx�ei�:Uψ0w��?@i���D_�Њc�aHq͵{|s#�XzhD��d�q@�+Җ�S&Z����7���	�+����K��R-�N�pҀ�q�J"]�rG%�`��rz�c�;̦@�4`�^��,��U�����a�8�	��Y߾x��nh$VG����P)U�	RFYn=�7�Z�.h�.����V�E�s�N�e��	�Qύ/M=����H�����޳ו��x�n7��O��[9xR�VG��⦧

h{O�H�$0@��ǟ���Q�N�1�t�5AH̲�/��߷�-[� ��P�T2�1 y#��z��$�~�\�>e����)��K?�R[���$�N�9�ȡ���9Bk�z$k=�{����<e���wں����(2Y�{�*|��t��&��%iX��R@��|eծ�<R�,U}W��#^��tMVǘ���R�.B�}�]���,��*1�n��QOܚ�Q�EB	g�M
Y09�<�|�n��'�.:pY��v�~߰��J����(������YeUٛ����������]�����r8��D��6��X�S�JAH|�X�f��j��v�>r��
ܚ�듪9wXV;w�b�c5�����+�>b${��fr
�P:����t����cV��!C��|〉`�13�uK�	>Zo�3�rh��8�����.�X��Tկ�́�=LLA�N$���f�C`���_��_^p&y�`#^��2t���{3�^�%�E��A��`/���6�����)����-d�A���wSp���*��>���������
�_/G�Pu'~"u�Q�<�E����\���',�4t�@>�e����@B���7�i+��FH�W���h`���])�#	�SA��+�U���������[8��;~(G����W({o?�H%\RGZx����Z���Զ��e���1�d�Q#5����l�N�c��T���$��dg���RH��E�޴m�n'zX|�E���/����P����D��cK}�x�b��*�7�Tg��lg�ھ����߿�y��+�h+��3�g���:���6�>v!+����e�y���o�l�?�»�Z]�Ε�L��,7��w���ϕ��O0�&{����ZeC�&���Ծ��\K��h8�I4�]Ydp�WB��ef�{Ь�TKoPnh~[�V/�\a�l&�ݽ�S�F��hL�_���0�w��8^(P�kBLO�J[�s\����)�v� J�d.���7%FDV���'[8.��ym`�T�<:H_)Q2�p�e��c��_�?��~�T
��s ��68P�N3ؙR}�I��k<�ѵ���V�(���#e<О�[�߮��2�>ES���<o��m� ĭ�@DhHSC���^������,�~�N�$9[mA�g���<�G^��	��v�4��G��6i��h�%S�%����Y,c� !�F�h�����uAw���?�I�C��A��B-.2��-�,�E�S�	�����=�
�t�#�Oj�S��3�3�,n�$�\pŊRз�׺��d�]�mvƦ�v������1����v��{T����z�A`{\�gy�u��	T���Г��y�~b!����z��Ѷʌ	��3��ot�_n� kO���6_�D�B9Of ~ԍ~I����w����2U�3�r��!����&(f7ۯp�8�܋P�c+�m��*xA�ǆ��k��gGPg�4��T�:5I�Y���v� F�<�ؓ��dq��-S�N��Fܺ��i�-,j�Z�ֳg�G6�
�Q�Q#쟉��-�rlUά��8T.��|?!�U�����Nz�x�WВ��L��m�ZM=*�Cml`tگx��+�8n���i��C
�尷���@�U��W�[
�9��)ޠ9�u��q��-T���I��|�{rn�Ϫ,�_�[{������vB�d�Dx��X[�z,��߀�y���M�L�?
Xa�㍫�T�kמ���C�5��E[K	ڶL!xM���� ]�ȣuY~����P5whzE��?䨅�H =����̣`G�O�>�R5b��ɡ�Ajxae�����ޫ��3٧�pg�N /�;�%���k/�tW
Ƈ$�'A���ٗ��LM����T�i��rg�<`���w�!T�����\+��x�ٗm1D2	T�Hz�emw��� n]�к���zeUe0�l����+�����D���Jmz�(#�e�����{��;����"�_y�
K��g�gbd���Î��� �c�r=>F*'$����*֡U�j_��!�^[b<�a�c��Ɖ� ���ݰ��jĈ�0q[5J��������㊂�Q��Tސ
��0$����?�x��5.B;=�8#-�"��C��c��\G�,�uP=4����/"xA}�������~_���9�H� 'Uey��^���ߚ�}�O�:��05��7&��}Y�����݉2�k�����y�ߴ�;���O1hD�����r�lTnO¬��4{� ���Z�j��>�g�'���(
i�ᰬS�C�8@�Ն*ݎ����b�e�i��M%z��Ǿ��� V�C���ܐ��pP�hFVj(�ܝ<�&��m��4&U4f�)ü,Ą��aҭ�oUk2��0Zo^����V���Z�Z'uBB��7�U�{Bc�F�.'2��';s���/2��s.4�GX�c�����Z��>�:��u
�Dj@����(�#=pT��e �jx�o���	]𺒆� �i' J�1GA�\�-���%?������uM�Ɯ�zh#�#YZ��D�m�� J����&���#��7	u��B7����������ܭ�/�1�^�x '�ߩ�9�f��3RH$���xy-]9��벅-	k���i8��/��z0���pڮ����½~��ǣ�u�lS���~r�U����QAF�7>�4.k�q[]/��/��������0��$���a���	��m+�m�z~X��=:gj���)�|h)�UC�`��S��B�|_}��RC̘<_�=�\v�U�ŧ�UQ�Y]����8�}݌4l�'�L�ɻ²�wu�|�m�HA�a��BW��Ⱦ��>�ۅܷ�P�]�Dh'O1ef��k	����9zIyL�τ�&�HUq�Pu�7Uk�N�9��g2}ω�Ҳ�o�1|	� ����������1�:��z�k��K�{[�4CDz�����8kÑ[gX&Aຐ_��&��4��=з��hx�qi�x��F՞�i�vR�v)6�â���qy�o�sU�ρ���ίJ��",�U���X�E���Z���t�@ ى���:����e��X����ݾog8�	ñۈ�J��+.V���s�[�p�ܠ�ou�� A�O�w�F�����Pv�K�-�l�/��\�".y�ojr
|��V���h�2�<aX�$�����f��]G���}�����"3`��F��:ْ�ôjv�j�)Xuv]�/���OoEɉ;����������}Ϊ�]S���Ý��$�%q�^G��2�������DTl̡eD<? ��},��:�<C�Hx������s[ک�:�:��FBYV���֧�cO���訵�p����Y����-N7X��!Z={��{9�*��(Eٳ��,快B+���|[5n���!;�$�r��\姏���DB5?Y&�^d�P
�]XC�b:n?	�����Q}3_��i>�8�f�M��z��UF ��p��C�Je�é����yP։xQ�J�����5��SY<u�<ʒk�dQ�9�bl�)�)-��7�7i6b~]��"PH���,��21���7���bCXR1�)�Í�Ac%�K	B�ԕ%W0*+I�F�5~[W۶`9�������2�"}/t=��n�f�2�N�֖#���(��n/��67y@Ts*,��T�3`[��o��l�Sf��:xCLw�:��+X�?�4�zP�Bm_��p,7�R�_Y �����f�"P2-
6�v0p|R������.I�)Զ�KUP쳸t�M�Q��Ũ�U!M��O��$�k���(S&ۄ�ce�Q����,i�ۓ-X̌�g,n\�u�'���4&��p�x�b~Q��&�u�xi�#�f�'ߩD^ ȀZ}�`QH,�����;��x��AU ��32�O5�O..�ǖ�l`�7��-'���j?Hy0�L����a7������nMl%�?\�,[��������jZ>ӓKr�uc���4�d�?ir��[I/z!���_D�L~{�jO��� ���\�
�����>9A����F��F�Z�`D�h<㒈M�"�`ͼ=�"s�0u2͟g]AI����$ި5���VFނ�ZPM垤*ߒ��V�Z6��pI���1T0������#�'laκH	��n,�m���$^b�3��"�*a8E����}��lp��2�����/>�u���)���^K����b�B�{Q�|����K��\�l+������+��������,���d9 p:r���it.��߀�~���%�f@dD����$%��a}�M2j��>�]6�`k��lfT��'�C���o-hp}���0�4��6W���A�]�٫W��
"��|�,�w��W�$.x	>��������5�� ��]BU��s���b@ �Oow�Q��Kj���5����I~�������ܝ�	64Ѕy8$/UB�����'_��K7��"��i$ҹ�"��)ɶ#�:�٦��UE!��`�3�MVl����Ŗej]ےoU�"� iViCOcR��^��7��fjD���sN&��	Q:�+�� -�TJ*%`H�����R�p�|�����Q���?�+��[��>���j��W`ş@��#�T�ďg�l�j>�}#���b7?z��S��A��Մ��߃oߙF�QG�cWc�seܪ;�&!K�����p����L6~p۸��R0h���ͪV�ե/�M��T �~�/Μ���>̘N)��@D����$>�y��!�6��<T���-˓ķ�Eagu�N�͢��P����)�}���+l�(V)�ɴ�Т ����zo1lx>!��`5�ut��Y�Z';��?�?��㷁x��:t��n���ף��^���Jeg���^���hk�i��4IFbf���k�}k�_�(,W�Na�&Oc�d_W^Q!t��&_)?7��԰q�F��~U:{�i�~b�^*�C1�P��h��A?�[�@��,�+lE��%�O)������S���*���~�+�ֱG�`��FҦ8����;C�ٶ;�#i!{��D�w���B�-3wcHvn������Q,��\#C�����҃��納���Fx���0n�\uu�~�o�\�r�A.�����SB!-U'�B/�ͳHX��7�h����� g�(�>[G�q��a2 �J�5Р��y�A{��FF�	h���5�+����mWT�����&A��v@����m���.H��S\�WwNM���@-�2����r��r�i�M��"��_Q�\fj��);ܑ�|�LN�i�Ԗ�x2�Vj�U�SV}� �)1�$����ld��!���Wni������v_�q�-02Bj#�� ִ����i��H�����߸W��gCLG���$&[�����U\�<I9Wi`�����^;��#����-|��B���� �2�j´�������jVm���޸*��F������NV1��bH9����n��0\2h��*�wY��nA�J	�7P{�A���k#�p��v�p"s�2��;+O�X�[ƖC�A!I�`��G���������
	}���A?Ee�V�u1��wx���a��Gih�K������M6~O����Q~�Ύ�揞����'�Rzά%�?:����^^�n�sU6�[Mp[�d6����s��:#��~��+$	���rr��d�����U�𴈺���}2�U����9�r�'o�=0M���� �Kt$�8Ƚ�@�A�~�Ȩ�݆"@v{R1��qsK~]�W��U��q|�3-/��p�-jʲ��f��؜Ћ�|�]��m	���E��*�Uʡ�����
�X�vM�ɚ��ֿV��ks)c#:��{{_�o0�8�]����uFY��K��ɇG�,M��ʂ%�s�R>�m��;=>sR.旕5�X��\̟%��QX�JF�� �fk�����c;�w���ZLs,kn�T��}�M��e8me��5�*�SƷ��$���'E}R���栙!�����
 ƈ샏�8�ȿ���З�Ϸ�{"b" 
��]e��'���Yn��� �L���92�o�V�Un�t�,�cG�D��ꄬ�dH)[\X���#e�o�k�
�7!�Ŭ=��6DAao S������������Y�� \REGj��C��׻�%U����G����h�_o�T*���I���c�4��Ӭ���J�zy)-����7�l��Q\@����<��K���c�[]�孹|BʓL��a��͋�ӌWɋ{�����R+B0>X�6n�s��V���b�w���;��Ƙ���<���]�jI�1 ���H�BL=_���L�(f��n_~b���b���p�|���8?nQ�3��!��_{�D�<��˅��Tք���t�D�6�]K�("F�>q���%P?�����u<+r]�bu�ą[OpLT�B;/G;V� S"�ߜ�x��IE��k�X���٫��;4�MJ�'�W=��͜[���h?H���k��/Z(�E%�;��F�d��O�T��PaI�RL40sPjOC�KGGߵ� '�O���P�:�w4N�*T�;~��� �i>��'
�]�.�Ͱǜ�����ս����a�ޡ�}�Α[��ç�#$+��ḽ��-I�_K;ˈ\W`&&���yU%ӳ|8ܦP}j��ʕ*��������w�@��+l���ɓ6�#d��&�~��L�xړ4'��z�O�G��їok�i?v�s�T�̀�v�B	���Kwϗ�|���jA'�tԑ�h�U��m�^Ԕ{{yL�'�T���PXOԔT�K�45.����o���%�A\��z�el㿜���*�w���[~؄���������zm��zP�}������"* �VTad6 v;l��I�N,9&��ܗ��Z�`�%R�QXfe7����j�ԱhA�E|z���[�m�O��ͯ������M�b�L�AP�������Lb��nc�-`U3�:5ܐ�}�b2�	�������1O)��D�ʎF�g՚^@4�9M�u� ��rgM�[��J'k}������b��_UMK�������3��m�}�%`/yr�nJ����1����.��5�Sx����e�i8��q�'��ѤNT����ݬ�R�A�����퟽ 7�Q�!��*�VK剆U�B��n�ո8��K_���?�%���<��O����K$m�`�HG�`��-��=�S\ /�/]�X�6��R��BL5���j�v�7Ab����'qH*<�8I��s���\hrnQڦ�RA�2�4�����Lǀ��/Mh������}�qSr]ayդ�	T1����!;�S�F��0��9�̌J?�����M VC�t8x�ؘ��Vzӑ�V���P�y�ę�~V��� �ٱ@z�V����z	�b�rN��IP���� ��Z�^!?�nʡsL#2Y��!Ӹ<�[�6��vO�BǟI�Q��ǓФW�p�0�!�6-���TS�[t��0yjֲ��#����V�F(�������z'Z��=Ԣ�a��Vκ���&��Tl�ٸV�@�O]������z�f���.��
�qU�[��dX��z�����5��;����u�[~=�����kB�����x��6�#O��A�D���Z��;h���S��mXy�,J��z���j�/a�����? [�:��vRM5�E��q��?�usf!nZ���W��pstv�"m���ޞj�e5�#��0K���&ӝ��V��>6a'�*j�p8`�Y�����rjN�O�̳�K�J���9#3OPhߙ5�#��PO*}�;Z�k��=M��A)�J'��:��?5�&z>�����0��lK���\i��꼔��_��󙤄�ie�[6W-�-RF��,�,>�ْ��u����	�x��ޏ�\��M�I���}�ro��po��	�ml��:���o� ���v����À�RH	���?��X;P�퍩֟�َO��w�K������!�MB%R�F2n�o�*i�-y�Yv%&5(L��CuZ�b���4��`O�oj�x0i)aVw�m�����,{y��խ�a�|5uC3��@������<mw�Z��2�jqnI�S+YW�H�P[����-Ĥ�]�K�*Q����&��>���F"ti~�
�@.��S\$,g��S	���	�%,�W��F�[���G.�4�x�D�B�P��=�i��S�=*/��!�b��g2�_���ʨ90?1�\"��i:�\|%�� ,8kvn�_�W!�LE��_\�U��Tu��ҍ���T�]��$�t��>���n�r�&��R�Oq\-�U����?��c�G -�˺7uʰ=�����^��Q?i>��:@�����Jx���F���8�|S6���h&U��x�rJ֎�u�ɤ̓s�}���=�h��C�x�M#��͋z�5�FzF;@9�W��D"��IN�����e�Ϟ��?�_�Lbܴ���G�e� �ct_RcĤ�t�����<�t.�f�\�8���<���%���F� G]b*!� 5I��a�����C����{!�xx�XM�=M�;����|�����Dk�v�N��' ��xh.��I��9=7�t}���ՌID���1|gݘ⒤FQzD���w:qL'�
@G�������ԇ�R X��<=����.�CK�bg�	�Ũ�W$	�����ιLt{�s���g�͆���[�'��9��?�������y��'�:��L���MȎ�Mb��b�~od���}s8R(7���士�PKHy�{�j�o� �g�]]Xv��Wݷ���J6ܫF�en;�Op=�.`v���
ͤf�0�M��-��������>P̟���4J m3�Ý��"�ډ}��G�d���e��?b��4�Jc�!l�1��-�`�䥱B�������Xys�|;v8�̵9Oۂ��,� ��/��_���%]T���#�HF4�0�������AN���%�{+�*�8ᢺ��n|c0TQ��=�U�@��z\���c��X�&r���U�D<;r1�x*�����%ʈ�k��ڡE�v*|���0F��0D/����V��B#�n9ܘR-�l����?.N�nm�L��lQ5I
��ѣq �F�˱8�^M!�HZB�P�s*$�0�vt�Giw���}.7H���Z:�DK`>���n⭃�/�P�:���� Փ\i}"���]>���AG�^9�mk-�y}�uH��|I]|G�.څ�cޗ��+X�&�w'��,�Y3�d���Yz����w�ׅN9���|u�Å�d���%P��^�.ѩ��՛=�o&#fK�v������V���f�|DxTO�r���w�wPY}v	��f}N�L��<�~�-�������E_��zۈJ��f�˹�3xg��0�b!��		*¥Z�YF�� �O�e_��87�`�\�D�c��+۶��=�J�k��$%�ֲ�Q��\Ü��C�q؊o��m\�S��~@Y�h~������n��<�n�y���^v	��j.����rh�"@D�r�֠~�����N$�q~�0<�ի�k��q~���kgD7������vs/E��].��͂��J�!�6�Wi�ׁ'�!�ِ[||#O�Z�<5�l��W �����]t�jR�Mm�
2�$���[�{d.���6�>tR]}���hn�0���^Z<�h�)�X�*%�W��b
M���;���e���3�Ɓ���:��X�Xh�R�Pc��9��G ���&I�l{�cN�{�[�g�"|ptW0��<eo7�m�,;���!��5�x�I���Q�����+U�H�Tz���i�~%��,��U�h�p�pa>��EJE+�Zb,�G�1ȕ!*;�*\ᝀe��������-\ߪ����M<����aeA�D��	���_i���_X:)F�Ǹ��l��+��4�IU0BE-v�E'���!�gw��	�MCvh�Ė���K�b7�w&C��� X6=j�iJ��u8G�j��Y� CT��2��8����U�1�W��A'ȍ˟N� �*�[;;���B����-i�	
�~�>fH������Y5nK$+:����o�5��t�R*��G+9���F-I>��Fo��Dټ��̬����*�΍ob�
�뼌�tO�j>Nݢ/i?YǰĚ[�A\�j���ǍN�W�j�%p��1Y'u	��}h��� D�ο��"C$�m�7))yЁ��G��(�����q������<���`�\�0{�h`|L�Z�g��OFj�,ٵ?O�H���4&s��J2$)���1.���_�"�$��j�|�X���F+����8�Ud~�`�vvO�n���.������Hx�U�]���M��k��_/�|�
<�f�/����i�;��ѹ��?׃l4�h�AA�X-π`��@��74ͬOQ��'ïyi�x�(��	~
�\���l��I08)�xՈ�?y��ϡ�9�Ӳ�k�;�p��- ˳�y;yS��4��aƊ/w�KH=���ڵ�g�%"�{���۞��b���/�|��,Ů��K��V��l:�pL�] U��\��+<Iv�v�T>5��Ds ���.�i�`�'cІ [��6 �v�O���H2y����@�QG�
���m�Z�ٌ�f}���Ǐ����L��G��,���	
��`M�}q�3�����Ѝ��?W �h�Q@�cf��A�jH:���3���,�]s�(|6�/�t�/�yZ5M�`R�A_���}�h��&�b{��}��1̗;#}haP
\�W8�
i��&n�7{(I�ݢ�Ym��5M(�cbs��I�ו��MB�ǻ�'�]��3�����S�DC֬ώ��sl��)��ɵ@Wڎ ��tm�2
~�bm?�S���i},��C����n���!�,ɑ���E��='�oN"�KVG�`o
�B�Q0��HxXۍl*�ō��%���-a�po�Z{�f"����
��vr��-�,Y�S
�1�r��]U�$b60����,x��^O�6��$�:��;4Q�"��4�1v�o�f$11��x0wp���bm�y*��N����@�@���KUoz�O���3��EŞO��﬩wWs8�&�n��K2�0���=\A��7P�+6=�=%�N!�v- �>�?f�" �'���)U�&�P�`�}/?�� 棜WU4�粀��hؕT���>k�����Vg����ƕ@x|�~��B(<Nb��K�����/�h��b�ϼA;>_���Pt���4{���4k��˴����
_D�$�;&e7���Վx+?e�!<�o�z��v�m<t�h��<l�-��i�~�q`���_D�{m�&*�� R��\�W���m�Q��g>��H��˃	�|,��4�$���|��n}���y�Q�g��ի�ۺ7ex��#�}�#���.G:��d\r"Ay���u�.�D��>5�<X�������.�u z���7�h,�[�OՉց�0	���\f\cF�r��FY���v5�W��a#�Ŷ�jӟ(ui��陼F���_�-&���E���R��̹nр�GC��	�JQ��ƺd8��J��w׷l1��b礑�\��ﲲޏH#��P��T��t�'���d�W$dq �y��-^���,�>�k����b>��Ű.B��:i���{��:L�_����L�X������8�z.�6�M��q�'v�]�󷠽`ɕ�����#]����NJ�d��|?Gz]4��C���TH��Ln�w8��r�+��U�O4N�(=�XDۂ�[�y7��b��,ײY�§mI�������_�Ӯm���l*)(O�+n�����1H��8;��#�b����5Cfi�E��J�+����=�s�Nղ�X�Jd���([#�<�90��8��7�V}�ޜe��	F'�6 S���;�{tR��M	>��D���V�����u�-�����s6y��{|N��Y���	/�����ɂ}�TB�,������c��;���#�����ܧ���� ���1TYw�w��nEn�4s�s��DLM�߫�|�k�4�M�\�ٴ	Y`Kf:ړ��)"���:�o�#�;r��:~���r�9�X�By���K���A���ȟȣ �̵�c%T��٭��_�T�0�H��s�R�G�uú޾>���@�*��H��{�G���&���� 4��{��B�ү���`?�GJ�� �L�g�?U�!Y���K�!���"=�C�s�j�?'ct�g1D+I��g�_��V��������=%Ս�L#�ed)6L�`������p]ʫ]� ���\SНhV�v�(+"$��R�G|��k��?���/GƱ̴�̱��7���uH����_>��\���\#p��uŰ�N8�;XEF5:�LCv��=��=9X��>ӱ|��݈|C8��_r��'��-�ύ���I*���5��SdV�f"�2���u��~O�ӡ/wTf�*���ߧ_Fb;����;l,����&�����BH�o���-�C�x����q��X�������@9���w�W�E�E��ed����'��W���C�iu>��Y�����?�<� G�0��v�Q76�)�A����3�̒"�ܩO�ʥ�Z�XZu@�Qa�X�S�O^A�O���Ņ�sf�޽C�l�����.�/��E(��0[���6:�����0bcu�3z~��e|�b,XB]���=�}�bR��$$f����D͎�K�T̜���v��L)'�^��2��sT_%*:��OE��̂�`r<�x<OB��|+л
8��:�X�rzf��5!g7�ac0?Z�:'ns��r?�i���}-1�Cj_w����6�U�-}e����1q��ڤ~�I�W�<1m@��N��ɉ�"�Y�Y� W�(��ni��
.�Ͷ����o�x��b*o��!BD0e���=�PB5���l(�� �[sW���D�gf+�)����K�h�u�����v���o'm�� Q��_9
'�0��� �x��ǈ� 9�eV�f;)�g����I��e'*fR�J`rqArQ�3�{H����:yz�r��<Ju�߃����k?��(�Mn�R?ry�(�'��]UU H�J��^JS>������cBO��n|���k
����c�ɳ]���u�q�U˩,��7�;Uwi~`�1��ĸ*_G�C�ä՟.HcAN4?�b�G�]6}>^��`"SWf��Dr+�Nȟf�����-=�2�n����#C�9�'Db���T��7gŦ�k��y�MO���	��~3��}�A��&���;�\QW��A1C����+�G��Kq*EX�[D׆|��Y��۠�	E������R�F�9�H�獪;�sq��k�>W܆;#w�@4�� ��O=覐�Np<'RU4P�k�YYs5�,��sW�<�/�JL�)���!ȃ��9-���k����8.�g[p��:���k��m�@�y��R�%��2��l�(��d��Xą�g~� N͠K�#1Q�7M��.�]���]�� :f>��J6�N��ٓ$� �z_�g���r��0c��$&�j-��:�r��3 �i�5�F��ĩ��iH<�؋Y�,�4sg�2�λ+�&�w�])6L>�R�{�,HNOf����3|����Qˠ���A�r�`B>�< ���$�y׌53��%5ȯ�}�g�mz���,6�W�i�8�Fbr��O�`��,ü�{)��y�BT�vnmI1W�t��x����_z�4���(�)SKM �=���b�摃���7�.Nݢ���x�Ug[�0* R�t�k�B�nå�Y���T'� )��D�0\s�_�;d�vBU�,�u���n�
�Z��&k9�p�DA�-��`�&��~�`�G�� ��z���B>b���3ra�����D���>\�y�Y����7����0����`
�k��������� ;�4*c�I}J�e0�&���io�B��2�.�j�T���H��e����!���XQ�r5B_}�{}6k��+��s!ڲ��J�8}|]A��/aK���.��C�|��еn�U�@L"����++���<>B^�^ o��@�|�K��g�µ�2��0�K�R-u�9�|��G�����i�徘��6u
��e���6dژ����Y+}(��߯,��Y���/��Dy�2񷀡J��]�挴�S�sK��1x�`���#d�S5<N J-����\��9��ٰ#�`KR��-S-k�fi��P�M�z�}l��h:��/돿Տ?�4Σ�a�z���<�|��]P�� #P�����D����WH^�'T�a0�Of��tV��|p#~>�Dn��+!s=���3 �)׿�8X)
&32]�W{�	�
=M�3ad��~q�����n�7���ie��N�T	�!�b%ÍNy1���L>Q;r{�DIlG�w�G�|� �T�l��f�+.�������, ޜ�;�dFr&�O�!��jRxNW�#�`�ܤ��֪���9��]<��B�F)�
�t��o�E���a�m�%���Zu���J~�u��V���7���L"�gW��zF�bC�ά2�O���ܾɪ@s�l_�ތ$�_?]�7��j4��c�!��_C��1���l���D��2X'a-����λ� �]�������挒hR���M^�ܱ��%�g�M}�լ��|sf8wH������w�vTH+���`ʖi%��w2���Z���$�@I��ԀY����4+�@�J|z�T�����{�])'ݶ���9j���T�(q��c�&�A��X�ދ͏Җ,�B���{Y[�c͕��B?���o�[]�7W~�%��S�9��l;���m ⷶ'���R��vM�����'D�J����ǲ�Í�0Ȳ��o�v���"M��ꀏ��}d�݆L�T��)�t� z�x�*���+�mɣ�5��콋�F�uB��c�n��>#��~�/�����$���ы.��%��h��ns���0+RE��u)��w�x�ݦ�g'���~
�D�2e�HW5]	�ؔ��Jԅ�B!As�vtߐ��D�������>Z�v�	m��O��]����sތ]ξ���O2fݸ�LJ�-�|}d�����kחՊ��fa��}.b��mn����.���W��q꽰"{DA���S?���u�uQ��I~��	��lp�T�ش`�������Lc�u!\~���9�܉.r��SsF
��?O*jL(�f�����v�,un&b���N֊���eԗe\�58ū����AX?�
���Q�@�}�t�SC#�Y�HE�`VN�k��mQ.Ri��絝�6�R�ŭ���T�c=�>@?t]#,:�c�!��"b���\(���9��7�Ӵ	�f<k��|�-s������Ҥ��i��Ǹ����5O��:�u����V�N��p�RĂ�O�t˷��W����^��8zo��_
H��寃H���^���A�&����>�u4EZXf������.��kP*S�F������Z�^U��nz���Q�px{'m�q�R��;��|=�W�!�l�K�
�쮸D@��{L�9�~�US�M�1��|�[��<弪E����=#�m Lk�j�<��BpJB�aݣ��&��;8��g��vd z�H�#�퀄�ݚ�Co �{�H��������G�_'`�R'"��/����K���s*]�F
J�?ψ�M�7�hwZH���m�^��CΆ��Uޖ�����P/��Qt7���/jjs<H��d~u5+F(��,'p��?�~��{���������<%��r's~�o.Ƅ��'�J�1�8�"���@�g��[ �SͶ��=�LZm��uV�a,��GY�DȮO�����|w[�e)�k�@�?O;��������~�[�5���#��,���/�J����9c{.V>�O1n2'
��;t_���b=�	>I��j�?ľ�`����H�������u*�FZ�F+Aę�8%��$�:�|���Ӟ7I�#�|�	�u�;1;ՓZ�80�vZK�����< �{X�f��a2��:.�W���YwYF�zdy��;邛�!��c��tJ�K���K��%I?��k�h���4W�~E>Q�?D����xt��{X�V�
���/m�Ԣ$�X�&c*���rhZ��l�#H�a�a��^�]iw����^/����j:HzC��P�ÿ�F��!r_��Z�ha���h��"픂�=��b|�h�qAf���u��c �1����˄��'�M��r��ޏ�*��6JU��l1�,Y��G���HT�}_��G:�q`kS_jz����O���u�vV�\�3o~�<b�W�{7��M%����[�.�<������|� �vn�R �L��+�:r`�b�\�듐m���y6|��Š��,������ 1�ɝ�cY#$�M���!2C��T2#pw��
.z��m1#����T����3�oX���(��9��C��%@BӠd�g�U��D7���q���˃�fg�+M�c �߫��_�?�b�x�����'7
ߴ�f��B��S���S򭊯�}!M~�Ԧ�ܿ<t^�/Z��0���<cS�l�4X���\���e�#R��v�a.��Wy,��|Z���T�C$�w	]A2-ۉ3ۓz�(�R�(3�$'M�|l���pk�!\�� �틦/z�|q5RD1��^&%�nSh>�J�H��0E��=!T�^S8��+�ײ����ru%e���^�7���?q����"���_����]��AM����� ���L D(��kĕ$�g��.v�dL��^~�ԜR�>�X׮Ĩ��Ly*+&*S��c��S�$j�)�NG�H�d������Mn⦀��[�Ps�BI@�`��R&�]l�ΡW����O��w�vӜ�po|Ƚz��g�]��ƗP� b�����6��g¯ȯ8!Y�y�u�vrI�T�A�(N��z�{[l�I~�$�kytJ_���ڶ*H�T�=�P��˩�m,��qd�y9]�,��)��7�RHy��ѸF��� �M�1.�~�^�2�R�w����=sEw=.�!"�/��sRR}WIk�>;��x���]"&
�#iO�M��Q���J�`c��Z�Ci�;�9���8�J��і��N��0�;���P����(��%�1�0�
u��$���]��x<�Gku�-8Q�J���3rfiu#��c�8[�T�r�����Y/�#�ԓ䎚"iׂ�o�3��$_<� ���Wͅ�7����F���	��Z�рt��^��!�䷜ojr�R�`2"�J��Я/y�8�Z͖qv;�z��A�
9pɞ��,��+��}s�^J���RgD-�ߏ�/��KWI�,����0�2���q��h@ճ4��+��p�͔�#)��^�3^��Қ�#�f&Xs��@�@�s��5�����'�c�|����j%M�5T�i���jW���|��G�B~n�x 6NԹ 01�uǪ� �*��|7߃���*n�j���d"��W�����f
*�l�Ûm������F��n�����u}����!	���`!X�)�`�3d��_��A���B��E���]�W?UN7�Z]���rdw5a����:u�E�mQ�z���U>��\b!���w6Ǎ�����_���'�˰y��=����1�ކ�1����d�Gt��u��TE�v�6��I�8mny�F���p��Dye�|�~�^mZ<\�ی��e{QY6@k�<�yF�7���A�0D2�yH�-1��A��բ�zmП�3��I�C2�cP���y�{�֝����]��L������fj��_:���k��n�إ�~��g�?�(~��nr4��)�����]<�����9T���>j�;߇T�ǫL��?�;�!��EN�`�s)[�i���c�4�5kf���9}>��٤Q��45?}ޗ���\� �s����#����w%�d���@0B��j+���*j��M����k�^1ٖ�l�O�m�\G��p1�Pܔm�
C�D�=�O�(�~��"��Eu�~ĵ�R
=�9���tu��/v��[���pZ�����gb�~w����!��J� � p(g�Ƃ���b��Y�MK%hd�r��D�7�(��M�Q-R��F	DV4��c��?���N�(�<��,�s8<�Nh�&�$�v-$E�9�r��`��H��Ѓ����	u5�a)�;��޳�����=��,�QQq��N�m�KiSpE�yM��T�$��8K�IU]�d�����(�A�`6�η<*X��۔��пt�ȹ��T[�	�!�Y^�2��ssB���fM��14y��h@�3}��'��ϰ�6;Ξ� b�{���5�-D�SV��U���T����Gp�,6���4��1ݘx�T�>[���V$��|����awH��	m9�h`ģ!�|�.ӛOd�l�:71� C�A�;7�J��v��O�;���ky�F���,�����&xğ1M��$d�\�@��;�I���)�[�q���D0xt��WKԢSF߯Jwk\�N:J(�y�R������Q�c�A��U>�)��U�;�?����Z��w���l�������ʽ�ѡ?x���%!7�9��o���/�=�8K�G����N�i�ܽ��Tr�����{V�)�)�㱡�"�ן�qn�$P�Z���}$7���xоɜJ�R��x~�Me$1x�~u/����"
Cu��ͱA�&�3Ǝz�&C�E���"�Vւ��M@��	p;�.���?2��_�q[��@��� ��Y�2v�A��ɱ��
%�4P~�iߎ��V��nӝBy�N��?���}�i"8{:2�&�hA���.UKʹ� ���[�%Y�җ먿��q�&��	��Vm2k��I��5)\���w �4
kj�` WO�Ҭ[ьtK8����`ԅ�2���9���{Rrtyz�W$B �9ƶę��+��hh�!�z���uunJT��,2��7�ȳ�� ��ݔ����U���|����;��_tkۘ�z@Z��ᓡI�b	E�Gcù�]�ĝl���`�����)T0�R �����T5�/É��_���z�Om̡�3�Y߲{�w ���l=�ڥ�;��o�c�X�(B�-�m��:�N�����8�)��?CdZ� X�ʂ�I2�K*h��˽!�Kj$|4U�W����*��=4�F:?�LQ���s�%j��!1-X�|������f��,z��:$�\B�3��$s.��f)՛�ꄦ��@�قR:�B-B�p�%�)�J^�L�X����A�[i�$�_�=�׃:�{�q����������&��EP��O�./G�����.SN_m��c�),��
ӎw����@tݕ-�V�éqB�iM�v��y�|�̀�B9�;2��g�t��ٷ�+tk[H?�ˤN�������D���$��m�
a�9��ꯂ/n�uʳ�r�_8��IkX@+��~�:��VP�����Kv?~����!6m�:%��]��
��_�:�.�,~��p��Ji,���S�Z�z���~-�{�
�ط��?�7�92f"'u���fķ��;lc��Q^�|R6��)��8N,����1(���A�kb�������R\�5���y鍧;��Ds@St�Q�u{�>}�*�Ht�u4��O��^lR��8�9j$VZ�prq�B(3�3:�}��x��#�MJ�4ѹ���O��3�ϐ>�W�\:Ipf�;�{�͈_�2lk�.��sB#�"�9�5���ӞT�-�E��;�|'4�<�5i/:	�8na��K���RZ$��V��
�g�ٖC�%A��>y}����6a���ƨ�b�r�!'-�`��	:�(H�7�3��mb~��`�h��7A��^z��mx�~�,G	�F��gN���a.
�R�܃d褞��ˈ|sn��e'��T*�U\�A��4�1�ut2(��Fn�t��1�Q�쀂x`sl��.!�)��wPJ���KV�S�&Ӧ��qs����XX�S/��}�����*�a~d��-���8V��@F�U�_<$�i�1F�1'I�q�g: �q�V� -��^�rߎv��l �եo�֍R����]�؂�>����zH�*N/[p�����{�M	/��u�s}&���H�Q�jYȁ� =��<��I���Mz��ZPz(���5�-�����B|U8�?�z�6(rXoG!!O��#�ev�4��(�U�`?��c���i_	�=4fq`1�ј���M3�1q�Vr��R��n�w�ԢԠOǟT0�B:�Ǒ� x|��Ls�ټT"n2���(��Y�@��1a�.k�	a���5���P���{���Dx�G\�hv���ǻ��v�[+�o��os���@;$D|��
�(��V�s<��xzM���Z и�j>�}|-�L��.Qoj#�����u��n�5��4�x!g�k� 4��N�C�]wW�qp���٫F�K����f�/�c���59p���/Rj?�P�l��ҝ�Zy�(td�=��]�8�Y�G%�3F�B�J{�	�%����'k�;i�vZ�8���� �8�?Q��P���2ҽ4�kM�c�l��)#�ʤ�.M���ͯ9&ƕ�4�@-\���)8G����%�:��ZVe���-�ݢl�Pm�^@H��Y#@d�]��T{��9f��Q�o2�M���r�%yZf�4��e�eT���Ԛ�)`|}�/��i��;!^�qN�Z'fq u�SLtIK�xk���Ľ�Q������?Ο	��a�LWA�h/s��t�q�A� �T� ���zcNZ+��L�}�ocRؽ�b7{5E��o�qt������9�#���7_���S���.2\�|R.޹;x8��nR��G��JD({��Ǣ�ӂ�A�}:P(�QK�<�s�9��X�M�U]X�sH.�z4�
��zد���{�Ms6���?��̗���U)��T'��������,}���v��Sx�rq����U:�vGYw����w�Bެ��̃��:������-y� 3��?0cctA�����H���G��&GѠ X�ς���]����<���gj����|�9
P�����`��<��t���գ�k�%�8c��G`�j�""#J"�c�o璭��ߕDoE��ŧ�wk���|�Z���g��X,�뙦��o�K��"�x�h���7`����%J�����R�Ĵ\y6��r��&l8H����(�Q�xZ�u6R���՜Lx��;]��	�� �@�Иu<"�sCU��q����(n;���@�xfQg�c����$I�J�R�cP�8r��F��|�rZ�)����\*Q�-���%�z��Mܱ����)h��dp�g��![:��g��J�%ut����yg]%�DO�0.H��l$�ux��C.Ц�뼃�*aq툙Q��*��3��d���R_���~i��nS()�y�!%�G�3 �I�E{�����RD��y���� ���IP���FY|�g֝dON�3:h�-�C�=�bV&A���+�4���)6p�&�XP����@h�C���'99d��ժ����_$��j��a�=����ا��.���\�uL���^���Q@��T�`2֮�A�e�uV>�{�ݡ��
��_B�P;^�2Ԟ�Tw��p+���h��%�l��y�0��O�pw���k^�.m��V�`�A�P!{�ψU!]x�k��E�G V����<pG[ީ���cB5x��`t��U�S��L+�v}������?7T��C��g$��o���R.F�x��+]�lw�z�|�s�����7�(�&��qק�� ��1F9j�qzrig�}k2��-�$���ߠtzy�O1G�����&/~A�Đ�@����&MCc���������~�&1�j���R:k#�U��=oY�a#{-���ӓE�\�i���lx ��%�kţ7#�"cw�\̈���@�;	��V���U6C=F0�]�1�X{�'�Fma�;����i�8�9�}�$�5��<�m�)P���!�;���5���du��,�M�!N���3U��������d��h�/���-+�7�[4�s���E��CJ�d��.G���^���ޛi�4!a���
vAP��s4�LJ�bAQJ��4;_�������7 n�(�4��{��B��vP��z�6o�k���߁0>�r���7R	��7o�T�M|�q��!s��?�<Ey
da"�<��{ٶG����z�k��+����WOF�#1�;,����'
m����-���JU+s��^u����PЛ:wK���#E��0o���.��D�EyOvO%��~"8��̗"}��`�����H���w���	/ډ#�F��M�L���(t�j��3��՚���I$G7#p~t����&'�ƹ�#�9d!?�K7؞�E�n9e�Xnyzb�{����Ű�0?П�W�Nh��ϭਢ�Fy�§��H�z���H��X�^��|��ʎR�*
���Tx��B�{�:T4��󶯔ΠHsCY��]��BL`��8������k�(Sy%}"ؕZ�jtb���Gj�z�$��&/6�'F��� �ꓗ��HnB�|�G��)��W�\�e�B3ܡ��J@��PUό���E�CF�\�i=A?hD�V���\*2���Px��7w<�ְ�k\�	B���ʜ� ���HBlp]�X,,ΊՎ� ���)"�jc A!�v}��8�FK`eS�(^��w��L�B��u��H�+�V7����o�h�i���_^��t�L��72-��Ӥ����*��#��f���/1)x���TEA�!��E�ru��o���LQ<-��Z���a��Ĉj��'A�icP]��ÎY�{��$��k�?�ص��`_e D�a`�^L�l�Ej�V|��T~����� lɷ=�$�$ٺSN�u��;>�	w2ꖧb�J�!�-���[��`L�55j&�%RZ�X$Ī��s��N�4fCyhh��Z��2V5�9w䒙��.�F��;o�*��jrC�$��f��}@kY 
��L�1� ��G�&&�,�a����W�+�P��~�����o��lQ�Z��/�0<�B��1;�����RRL=��RB���%|��`�ppK��2�\�����h� ���C/�oe���t ��q/�7#E,�1�W�W��Y�{l/q�dŕq�����[�_"MT�C�P�y�~����OYr6�Ő�\ŋ+kL�2_5��D�_�>}��Pf����2���Ѵh�E��~����\���z��nBt��!�Tn漣���M�v���D���N���39]4���括�5 b��9miE�{kpi!�W��b���E��l���<I�F}h?��EX�c�^�Ɵۺf��?�z��7)+��2k�su��f����o����Y7��6ٜ�Q�@z!�E�	tQ$稳��ڞ�뼶zm%�� ���E������v��Kg��<���ϖ�pz�'�W��%X7u#vg�
�M;ΐ�2�'X�Ԯ �<3�$�����cg�v���|2H�����h@?mW::����2\�`�A�7�ǶC����7� ģ�ztn��W_y�(n�B�\��ā�Di��H��hK;I����o�C{�m@-��6��S����2l-�%ɐ$M?�E��oe��h8n��Iv"����=�%oR1C�g�"NF��v�;R�TM�X\֒a�L0kF)��r��ZL��I�C\k�Gk@d�A�9{��H�M��$)l�W��ئ�68~ޱ�p��̕e]�oe�4۳ �����JG�rv.,�;�v尔��C����i��z@��[q<�N�@�ϑ��9�R�'�d]�.=u�f��Q�"��ڗ�8�H�x�%Z�(9F2N��[�y��S����N 0�z�����ݒ`�q�}q�eA��r[� �������dr�"ќ2��=f7i�	!��_�,/*���k5��8��L�l*�������T�o�����q�ފ������LpY�6I���_�o��7ު����`���}+RYs���
-�5��0��oId��H�+<	p���fL�ȻKn϶����\e̸���p�b?�k�?ߌ��S�����('�?p��́zh%鱮O�O��;aU�Nvɜ���Y����d��d��>�c:� ���Hs���h4��4o��7C(x�<G3�:$oy�1�x����938���	�x&X��``���
x�P��p�}�&�T9c�\�R��Ld+VO p��=�/�6��~?B�a�<+ � 5o�0�T�wV���y���k��ꀦ��`�j]��c���o(��k@:]V{~G����ڌVy!�2*�k�@bNT&u�N�Q΂Z�;o���[~"�=�%����z�	���^�O_�]	�>d��5c�2?^�o��R�L�j��=E  PN'w$��ru�n*Ǵ�Kh���<�G��K6�Lm���wpdӛpM��#W8&��i�#� Mw��r����>%(��>�/�?��T�g��>��V�)�/�࿴��n���]�v�@G/���N
�����a!��>�p�]����&{�����v����#��'q|`e�ֺ��ɋ'�Fh�K�@|s`���p1}� 6�����]YUX���:3��� `��%��18��t}h�|�j��suEtI���3�-D@�D	k]��j��o{�z`���/��Bm�	x�*��Y���_�T-�~�XB ����i0-���\�f1���&�]ak�ZoKsB�}_,���F�;p�p�����.E+$w���`d��Tc��i�N uA[y�p\������PnLzN^��M���u���jЌ����ù~���NUh��w��2��+��J�,墍�:1[�9�-Ȭ	YC�r�`6(R��Z6�ӚU�({�cuC�JE��7��0�S���D��-�� ~�n���@	�#�*���1��	{ǳ�K�;9qv��V���F��ERo�#T��,xD��(H:/�<�ޫ �72�%蓜?��@�f�1��RS��l�\E;�4;�^�3Q��vݢ�w�[���/�����<�ٓf0��^`�Чw�9�Ixl[1!ӻu�-[��Y"�(��6�ԛQaeɁ�C	2������P+(���nZr��A��ݿM;��}�ů �II�Y�p^M�g�D�i R���o��2m�ɲ�0���]��w?'���eM���U>ȁ0�R�=�A���{�@��n�:u��n*�.<���!�^Q�i=�-��A�>�	�z�u���W���i{/���Y<jy��k����B�ʪ:���b���VAt�N\�S��HꏚG��Vޘ�N����rF�����QG@H��[vu�����������0��}�"�V/�3�
V����ƪ�uj���7!�]rM�C�i�i.��Ir1� ��o��B��c�{sj_�絤qc��-�?�����d@�og�]����- ���2���l�Ο��ͿA�X�M\�sت������v�c������/]aׄ��f�櫅 ��!����snv HZ�@�k!dYS��-���K�-�ƃ0�H�S��ޛ�غ��oW������Iπ*��r8�<�:�WH�$��w;�+��b���n�sںF%���]�%-��{7T&�?�����k9�^�o7�g�ﰛ�֍��qO48�tt). �F2sn1pH�ֿ�hm��Zs̈́��>�gE#�!^SRt�b�l5S����=�j�^�_�[�"�U�s�t����ӟk6�C�� &^̘���i<,Mܲ�R����T',���\|bY�4���56hp���-���a���Z�w���t	��a^���M�Dn����w�.��OB�m�mA��}R���8M�"#����rg�j�W	�����')LD�\Eϟ��2�=��Ā�qx�I9p���F�a+/6�l�F۴�;��ر�K�\n�_[�5T�Ǚ��ʻ|I7I+��G�4
�4���/$J+qZ�E��)�";�����VqP8}q* �o���@��݃�:m�@SM��b6jX�Ȁ�(��p@�%k��a�jl�`�Ϻ���_�2.fk>�x�?���i�Y�����#{BG�E'�
-��2jt� $D�
?0�ĝ�E���O*1'���H3�3^�	/�ֿt��yN�&��k���g�L��_�$ԉl� �;�z�����p6bJ�vd�{�q���v��/�E�Ā&��č|�`��z��d���A�7�s�O���p�<o��w��`��#��܂�
��ʀ	#�Y�2 ��9��H4�N
bUR�1^�� �C&Ť��s�)��UX'4����ێ2dq���۝�62?Vi�-�i��g�qu���;O`+۝�2}�m���=�>�T��`�^8!`���Vt����W���RSk��|�9ɴ�'<�1аy4������7yイ����;�o�)n1�ڂ;��@���u�.�R`
)�]�E{�0�'=Iw��&�K����XA�>���Q�bz0Q��t�l���Y�\6�ȼ� �{���i僒y�_3k^^4�_�/a��c��5���%uE�8S7���lSE"����$=`��#�����N�Kvw*����,�@A�>�I1˖�y4�����N�@T&�� C�}���R��-�:�"�i�쭍S�O$��3��Ds��+	?��
QVa�+��y�G�pqΣ�p�ܻ��4���_�� ɇ�N"b�=W�bA&"�m�ϋ!W*o���=V�Z�[�K�۲`vL&�(}�uuV��<`讣ֽ��S*�tNF�.��H�X�j7$c?���F��>, �{_�]��a��V��3�h�{�>�8�]+��qt0�e��=�����%m�C�[��	�'9K��	0�������612e�����ɑ���	P9PB�Jv-��m�݋.[��9-��/K�LЎ����7�n_0kEP�[F�W�MhM��4�Ъ�:�������j}ޝ�7�, �0�{���顓cc�K܄���X6:�x�2fxŚ�`B�מ&R��~�fw���1���'��Y�-:tZ��ӭӉ���)�%����xYx����4���,�d�m5��e�����x�gM(+q��J J�3X��ʧ�搑�����V�N�s�ranu���nh��#�H���i�\���i�0Cۺ�G�:b(R|��¸����{ )T��=���Te���<�����T�-�0Ͱ��J�E�X7*R�ƛ�if��k��xi����h���l�m�Q�})��~��U�	���uG֠1�f���˂��U:��A]~����z��F����)�̑�{��|�E��*�8�o��=	@��e���0|��������)2�0b�w�����)��8�{.,VņPazJ���)d����;,����G ���-�x�jT��8��,�_t��z>mKB�p���eAD�Wd_t��m�8�n ��_�����f^�<��<�w�k����>G\J� �uF�`	27e��f�o�<�Xr[���]ye&QÕ�g-'�X�F�񼷢U�`w8׉l!HT��H��f��l���e�}�	4d��Z�;�;�����(����n�2 ��`���=���Һ��Ec�����ϝ��"}�����H�a���ls`�� j�l ?�`	�H�7��N�mZ�V��0�B���ӏX8�ي�Bв)�˓?������jp�X*��s���� .1ٚ�r"?Q��e��	Jj@�L�m��y�ڸ��Mc��&��$��X�������g���)�uy�Q<V�u��b����e���M]Ga�Ɔ�8s�T�P��ob���3m}�L�fݐ�:f3�o,�G(�X�:���k�k�P�<'��+h�g��ଚ&�>�����L��%����!����;�^^����.0�7j�#c!%l���,P������9�`��J���r�3�E9$�A��`<�kAV�H�9VĊ$J�J�����I�B)�A�>,���UU~�#\���i�,�\b�;n-^,x�p�6��*�����$L���rR�"S|>G���P�
5���ꬾSٹ�c$��I���m*KP�<w�ҡ�⠟RR�
8���z@�q��� B��z-��|��u�\�Ms��g��*�&��P�8+2d����%?:w����$�[��&w
�G�j�#�\[M@�,/k���ág�U�-�7��L���}��sK�[C[��<7W��l`�k��.͗[���QC���"k�ew�٦a���ss�^}!_T��Y�,��
��-ބx�Z0�c��捾�OP���M-�	��]��4��1���r�	���@A����w,�����������q����%�#�"7�X���(��d��O��A�e8zݙ�61�e��STZ��_KN�ۏ��W�J��8�/�2rH��{��> �'|G,1����]n5{87ڔb%)(|�5s��1��L��� �y	�T� ;0O߾�.�h癱L�76ғ�M�,#��0	�9�-�@����S�r�J�ݯާf����V�Ķ�u}nX�+���[��Z5��,;��>��w�.y�"P6N�1���y�(~�g�yЕMb/�aRn=�����ss��f'����o�ͩ�zA {#K5O~"�&�WqRU34��ʼ'�z���4��& ݻ�M�6�������A�;PJi�/�wET�'�ٵ,�c>��k�!�V���w��~�d�T:t�.[�Ƒ!^�{mCrƊl}of "�4��B�]�̻�o��x���\~��0V��[��ͱ��nR���rܝN`'�ޗ��l���&�#�_T�����<	�"�����1'���3Wn::Bܓ>�IO��kY�_Ȗ^1l*��['@ۀs���M�Ğ�P��0_��ۡ[�c	LO�%R���VPw� &�8b�d�0|�D��p�br�#��>I����az�?��	�_�/jr	�����,�}�v)���l�e���ߞ�v�_���
�J�+�եv��(۹C,�W*Q�,���g5W�7z+)����T���/]-�r���'�\��V�E+�'�<VO����W�2�י?~�`A�l� ���X�4N{�� ����6ψ�JeN�bGi��b6�U�Ƨ�I�MG�X)&z��uı��38���5j0739蝭�Bg�ߐ�&7�U���8���Q�hMF�s��$��z��g�����0�d�����PCq|w�^i$�d9���{�(� 	N�f!N�|�@�Xl�!�ۛ���D�%��"���D�R"��w
�l����s����n���b�>�
�V��Fwf��}��A�}ܩ���c�[�������������vמ�(��r`�-���0R��W�������������er8qt6���gc�������)&��M��/�5�sM[�r/�4Kk Y0ڞ?�\(��<�p��>�L��YwIiy+B��8-Zc��ڋ�|�h�B�(��{����>2Q�&��\�ڐk;�)Wi���"�Q�g��%jr�������f��ߑ��}P\  ��s�1�B�}F��D�+��h�}�F�-\��[q��b;%�G~����ƈ=��b�����M��-gw v'�ny�-�P�Q��Y<w}�'+zc�e�'�O�3|S'1����p�N}��{;�D�]��V�yJu#���B0���md����4.ER⏞
>��Au<�)��cx>�m��g�NB93GT|��S��I��	����h�1��$��Uu��'�s�U���	�K+xF�y.��0|�E�M�rO>�o 0�\>v�
��}���4"�f?�O�N��T�g�� �9��Յ��>����BZ���+I����ďW�~��Q.���5V��p�)�2���:�;��
�`q�H��q�nrl��E��	V��!|��"Z���kTH�g=�c��ik�Lq��<��Ȼx[�ގ׼X0A�j(4g�&u�\Rn�P���,#�5�y Ƴ|�)��p<XP���p�ިiYoR��~����U��zFT��x�qˋ����H���Y�z����R�#�t�_��Q�U��#B����������W^�3�R�z�zbV\@9��J*W�l�gB��N�o�wo�/@�PP�Ҁ�g6K��_���R�r��j����"3w�H���@��*:�l=i�5'z�1�(��$m�ء��e��[ָ�HH��1���Ϫ�����ĸ����vO�io�j!�z;1�.�&<�+����qyPY[��|�Ǽ�QH�_V�gkkw�Y>���3@Qj��6�%�0����/�>E�����g���v���R���g�C�G�E��3���������SJ��ê���r,�4��� �V��-���PR�n/y�ȥ���ݧ�B3�5�/Od=��D�u���i��� �׾[z�m�~L��q���mz?-�%깫����>����,�J�0bb c��<+��� ���V�U�9��E��g��é�x�5P����K�E��R�1�d��z˄%���p6�e1��&͌m���h/w�N�)W�����TP�5O���#V�Se����AX��l�b41�6���)ɶ�=8�d�+��:ޞ�_�ۿ6��OĂg��N�ϮZ�{K��܏A��j�W����@�,�禽1X��S�?�~U�x�b��ė�h��`�,;�z&�����Z�.���^��7v+�p��3&x��OUa�b�q�O�L�Dbj�� mf�t�,I�9e~/�S��K%v�����/�\��_T�'���W��%��uZ��C+́�-��&�g�� �:�TJ�s;�1��2(����Y{��XQk^D��"va
��LL�mc���b���Ʀ`�#��$%e�����B��c� ���!�{���h�pT_?	,��k�!�]掜�V�Z�͎�������(�q���e	_N�CX��� 3�di
��$�:]���gV�kJ���u�߅���Z�~���h����6���"M� ��R�U���?�<�?����>�a/�����u�d��)��w�9����6����q%���֦�U��`/I�fS��*_D3�A$�F��ۛ��	=s��H�d��UzѨo��\9Y�d� �I΂�m�֣VM��ٯƴ4�c��vC�Q^������d[	j.~K�d��ҏ�@��w2��&
��f�A$�ۆ�^wY���o]���P]�D�,���g�)w����	����EB:�L���*!�&5��C4��N��x�H[��&<�7
���q��A�߼��������nf����,���s��kcZǿ����%�'��l<�RY-�T�I]�T_?�{܀<b��Q�0ux�y��2S���Ҋ��3���p8��lT�'��o�g�Q��!Yw����v�����'kX���Ϛ�IŐy3�<��I��roX��ֲ
EP��*��p��GOo�V/�@�!^&���S�f���?xV;��s��$��ϸ=,�c/)svU#	�׮J��k���dm#�<2T�������2_$95S�ӔI>� S㾑jH1�K�˖�����'[�L�h�M�����q6U����K,=C����=|��)b����(UWU�qQ��d���ea$K?��)�&�p#u8�������`�˿��&ۄ�L��B�Gٹ��=dc��d-8^w�sKU�=�i~Gȃj��w�O���g:4x�`^�/�ϛ��ft{/�����&���۬� ���������d�a0�}��S�6�K�B`M愫�u`F�g�m%������6O����v�p�:����n�A�9�\Y�d��cZ.1X�1R/l0���Ĕ?<4�U�h����y�u�Jk�RU�5�ټ?�:�.+@%�.^�;t�I�����Na���[�`Q4����˼L�&�M��-���נA����ʚə�)��1�(��Z�C�kn�XWa��ΜN�-Zꝺ[�y�X�粁�<�G�)�/W,�E."��������� FW���걉����1�-5��w՘��#@ 5lJRfg�sdqd����v�G���/���,��&���L�PW,�',!qSg��d5N����[���1K�7�A0m@7U[��c�o�m `����@[� Sx��Lؼΐ^�e�W\.@{a�8GV�B-(�	YB���G�~٩�ZL�J��@��R�T�"�!2d�[����� �ꡘ��V^�J�I�Qӆ�.�.���%ZC+3
6ه�Y{m���|��0��P��q��:;��3�Sp{`��5��:���\>I6�i=��+ni�l�Q'O�@<_'}\.��1��|��re��as��)Lկ2C�iY�WnG~,	L��ct��b�8iʠ,��M)rֆ*4q��'�]L�<naz�֌fu2��c����[7�kEv�u�f�{��pl���0�F*z�g��]�D}xLɶ��0G@4ѣ� ���|_fm �\���}��Ŏ�I%�����n�Α@��7�q�Y�U��؊4-�4'HUM�iK�B)x�Ⱦ�����wjݤ��*0�ճ�T�)���,K<���f#� ��QxD>�Д�U>��T�yE)�����(�[{��DLT���=� \�X�M���>����=D�v.���k�!�:s��&����bw ���Tk+#��s���}OB��?+T��<j�Ly���H� �z�RB��)Kŷ.�>
���8=KI�c���,'/&ލ��#?�&�]k�O�ώ�W�-���{�8�E�� �t�r���<�DX�'�/�n,#Xӄ?���݋(F�JƦ`(r�W�ZN�;�ř%�M�9�ȿi���MI��j_�$��?��e/�{\�a?�"D���`��_:WE,Q5ja���km��tn�*�Αo�^k!��A�kb�YUn��:	S��Kw��ctX'��_�*<���Z��t]�ȣZ��+�T�w�T.�k��w��D��(���I<�Α���hZM�_!����5�Ec~E6������LW�KW����������	|��eS.M�l�*P��׍������02B��D鑦o%�5Ih����+�D��g0�� ����avT�:Ӂ41N�<��wy=�f��BB�^k�u�����j�|f)��'᜷��u�k(@p�>�״�
���$4�F���"� !���0���s츴�����e[w��ό�,-�.�p�|�
�����@��q�I�#�5!���{�������"l>_Ͷ�>������I��k{&���$�0i�8Ce���`��CZ�*��t�����Z l�@���4�č�\���۸ţThs�H�t��M�>�E��s���h��|��X[�w>� ��$Z��GD8���uKmY�=��pt.3���}m��o��L�s�qwѵ�}3*\�ö U���;:��j?cv�k��
�9<�ȡt��Qc��,�VfA�Wm�m��S�g�X{�G�7|����0\d�[�����R�ȐG����T,K�k����ރ�=J�!�~3�,V+�*�#��{Q��0 �|��:����ϖ���Ԍ�*����W��8��D?��6�?�i��v�KRݟx�Y�Fʰ�A�ST��3�B]P!����Ivy	����x�:��ɶ�;��y3�H�£ƯP^<�G��	ݻX�~\P���ݎ[�+$�;����p�Y'h�:�zv<����a����b���r��l/�I(�����/v��[�o^�(�_|8&O4�Mܢ")�_�:{�@�J���'^��;X���Uq��|���AL�I"`.9 �6��2��j��^��SE�x�0��01�L);K�@t늷�)^J���g�o�:@�c�F����ǹ��#�y��Io��S�)��},2}<&�݃tV�4�M��|.ȗ�k�j��pu������e�Z�c�Y3 ��C��<c�7�D��Oc��c|�'�ތm���1N�sp�=��9�>�NX�o0ӎk�f��ͨ�"�A-i_�y��jޛ	$WH�����'�4��f� n�7��P%�.ev�u���(�w����;5,~%T���1��8���;g*]o�|5��K2��68����6$L{���FryK��aA�����o��V����V3�4����u��vɯ������Y��B�oW�w8�9����]L�h�3��X���
�$��z��,�0������ȱ�d��������	0�҅�h���Q �b��M�����Ǜ岞lK�/K��/*֗�<�a�8.vch;<�a�^ͦP�C��2r�9�d���*�����Dc�f��8SȔ��n?��g����9��Vo(�yl~v��.\��V�����#�	���K�ᅙ����"���/��ahK�g���`ޯ�%����X̔W�b��b��%�E��߻%���O�.H�`7(�޾lԚ;�^2���y1��.�������"��!����/Ŭ���CE�X�YhU����
M����r��vN�YA?R���ʬ~�jG��POZ�u࿞�nP��x�R���?�xm~�\*�.d�ݍ���{���k��y�+]�U�߾Xp��GjfqWd(1!="9sj��C��l*}x��mr�]����[�4<��WWQ�.HD8�ޗ�A����yS��-�x�I����\��e"ߨ�L�M'�S[F�?�;m�l�l������\KS�0٩s��AFP#�j��3������G#�I��8��us�Ϡ�+��Q)(Z���8N����T�gq��\KSc�u�7>��O���g���\�����r�@gDu���|;X�0���^���h`H��������ԥ!�8Ã��ݔ�� 4(7R� $��ꪓ#��v�xJ�f��]�c�ݨ)
�O_�fu�e��W�U��ywP|w}2�nv:���p�Nm{R~ͷ)����n:Td������	؂�b����<�g���m��8c�x����w;�) zN�t�(g�n QMn���pmRg�$x��\)�)�̊�=��oő�%/W���O4�p���E }�U����p�/����7)����'��N����~�� ^נ���PU�lP��;q~�>�Af���* 嶖�a�)-���і􅤫 ��/�zFkwh�y�ׁ\tޏw�@����@�޲*�1��ڥ(�x|�_�"��+�P�B��Y�b�f�U��!:�I��ƹ�E_)-b��KwOc\v�R�'׻�����]R}V�G ?7$�^�0���_2�ڰ�]�,�^�
��m�_Q��6&����u=Ⲷ]��n�tعi$�s����%�x'3��a�!x���*!��v5N]c�Y�����g��`�ţ���&�{ס�%���()���,�O�<��8tB*�����K���.@��R|t�ːMh�R魓c�A6$����lH{ �Q�Mi1�O����Pʬ�C���$/5�dyU��M
U%A�2���6x�ȁh׻j>��J�3�&p?`�� (m��ٕ&��%x�;93���8Ԉ��c%C]��s�?�c����';��Ҹ��8�{'�r�4b{��째g����gQ��oް��{�;���ڮ!�8]�68��jDXrA5PC�|v�KB����%�*l��������C�0|�����<<�d
 F�N	z�M$5�� w&g3ÈK�^ųV��gsO��ț�P5�yH�8��~��V]�#˔��n�۴Hy&E��l�\��$�7Bµ�$�wr'�F��8���{|c�#o��� 汊;3�n��
�`�*5D�Á��Y�5>Mك����;J��v��~v3{}���}�%/���t9���&D+����"��Y0H�*�%g���z}0"���/ ]�����*�6B�0�+�I�M�o���Y1�c<(��5ی(�U�����m�P[R1h���IM%)s�_p�niz~W&��R=��94�B��̭�T�I6��x��� -�?Uu��+\��ݥ���1���I^{�D\e�HcT����F77�]��c�^A]����o4�}�����Yl�K��4����=�7^����~4�9U֐K��:�颕;v��*Up&L�Z�= u^"�ڎ��T�b�����w�|b��q�u�d����(Q?�J��3��_�-��e^������eFE�%��V���\�^����f��&fE�4yJR��B��/p�*���a�j�`!���^�aR���H�#j^���Ƿ��+����lY�Ӕ:�q�Z����	ӥ�+�Pu�ӄ�L.ܙ7uc�jC�T�D
�ک���k��vV��j��<=��M0�F��V�1���Uյ|f�
��<����7�����lopO����|$4���촷���N��F��O��ʛڤ�y��jɪ���4����o>��J�|z�*Q�����; �1�,03��n�S�L��y�Ր�T"H�?��)?|n;ݞ�b9��~�#4�l�7q����౸��O,bZ�|�re_/q��'Y~t��w�I>C�x.�������;MEF��-�	�����Ǡ���z j�5-�r*�a���]��{�ovb����	oep����R�f���3�7_�a� Q�*���T�ڑ�����X!x׊���u��UR��� ������K����5At�NLGo�,�|C�>u�D�G`��N���W��B�54{���[�b������Ƌ;>GJ�6��y��<$C]49!q�x����G-�]u�	�m*�#0��I��F�0��t�8�����#�lSP��7�¡��P�}ldR�����*�K{4k� M��$Ms�["gHp?����������K����W�UT���1�������#��Uξ�r�2����JS�⌎)-�QDM�J���f�=����W����AB%CSL�J#�U7~��*9$-|�Cz!H�d7 �D2X���Gj%&Zѭ�\oRG4u�C�����a�m��T�+J��:)^)ભ� �]?O��F��Y������}�Ǎ�����T��Ȍ�N�W�rّ�^��$��V0�$f�1��d�͈�t��0%E��dzC�l�H�B�P��'+U�h�C9���D������|�Ft���V�Q3��Ai�x��ٟ�*��
H�AK��� ������]F1mݵ�%�L����a��,�@�����#�U��%�sU�(x �F�q��K��R� �$��y�9""��w_}bR��3��W����ݾ�Uy���O����7�9��-��ebhS0e�XR�C"=���ښ>B�:}�Gۑ��m?Ħ��Z?�Z��`&+N��J� �>竻[�9���:�i�X�2�Bn�!�L?�Q僘1�Ϝ�&F����]�釳L��:`���/�H��K]���4$~f��Z黕��� De�e+ZT���J�~2�i裇�i�˪�⡏�2As��v����,(N��:R�Ί�
W��c=��hp$�Q��kGn/N�ur��|0��=G�ɽ�s�I�>;,|�H�L����vյ7�f�F�2ݤ�	n��eJ}X�[1i��6��Et#�6\����t5����ܦz���)9>���{+	��L�nM�5Ѯ�����!�|�j�ܔ¦�43��,�x- 1!��%{�.�ј�(�RJ��
�(t	�?8�2��a� �,����%<�H����g0QA��;�=Ȇ�h��=����~�Z���F���#���e*��8g��$�|^�WT�a��ɷ����d���u8��u�/��K�I������^��09��h���E�cb
���\S�K�f�!��A��|7�M?�6�p8�P@�hc�h" ���.�~��J�7��M���6��?�A��%��O_��Fc<ӕc�c�
�ڧ|���r��L��8���E��+7�p��'yTy�2��{�Vr��F�Q�m�����ˏ��_5�I����־��`�h2)�7r	��jA��t�p��*� �^#�y9��d�ps���<����y���Z��Y�~�9��|�o��F����5uHn_e��}6�����z��)��`�_�ل<m��:X�T��e���B��UM��le��d혆�ONmᎌO5C��k�U
r�8��?��ߛ
?Vs��ܤ߮�p�]_X���F<tt%y4��2kpC丕&&+%�H�n�н��A�6���ޅ�u��
@�F����^��;��x��`hj���c���>I��е�gS���9�>C��b/�o�:�F�k�:�ٝ:0��\x0 �O�uFTx�VB�-?�Vi�4��=�_�Ǣ��J������s�:��6<&n#�#8�?/;J���+Z:5�;L�n��uYY@ej����0~�`�d����ovx�t�o�8��8X�aI��=`��f��Y�-�n��2�s4w��c���m�ӁQ�TDH)���Z���jOY�F�.c'�� �S��e^)��?RN-��[MBh�g�o&q�X�3�cci#��h����"����k���E	��q�Q����Fz�K4�3m���Y���>�����!�#_<Bz�O���Y�o�d+�e)y��ǧp��q%yRJ)��B����*<Ω4GQag���|/�m�%�U�����V�����0Rf��e��6N�IjC�KA-ظ��쿪��6�d���u�yK��G��W֦�����t���ч��|��R�h*X��^�8����Srw���������ؑ��	�b����~���A�B��1U[\�'ת=�$F����8Nն���������ջe��@g}�T3H;H��n��);�*d��� D�s��ܒ�"j�G����va�:�y�w±�����o�8�&ö41S\������"�5�� 1�ɢ[k�vV:�OĈ�
a�l���s%�7�xB��t��V'R>>h���D����c�]�*�5��n��\�D�K����O��\�s��y�)"p�_㓾��X��H�Հ5D&��]�>�5�NkM�b�A=k�G9��yn�L�w+�4�A}<��f[����hZ�?��&_\���@{эw����&r4j5�㑠��#c�$�,*�`b>�y��迍d6�Eg�&���C�]0�����C��+�4?�&�Љ��&b	�tej��m���g>���/�0�f�?#�^�����MkfĠP�<d��F�I�bL\G�l6.r����(!<�;��'�q�m����ᐲ:ou��� �6���;lT}�m-2�/�fK���OMb4'�B
I�ܫl���q�BJ�<	��+h�������4]=�Z�A�6�"�Z�6��c+@��U�54��m�nd��>�QȚ{Y����k:��\�����,5�J���������>�Pb���J)�s��)��1`���q�^��kM�u�%�7���RwT�P+�}��_�o��q�1k9���"dڮ��ZR����ś�DAC�C9�<��y��@	C$��c�聛`�(�rjy�=K��;:Z���_���\h̿&+H�Ծ�l�V|X%��#&���i	k~�e��I"�]`
�ָnR��. �/�����3,���O&ے�p�L0V�e��vn�̕_�_x����c?;5	��,ҵ�D�m%ȿ� ��sf ��M���f������+ߴ�7<z��g�i��������c����T���4�6�E��������SZ�qႮ�YP�y�LLCS����A�"eU ҁ�@�?�R�)�ѓ/��������(��>������G�;>���W1���lZk
��f~���t�t�5�E׹��)V��z������.Ź��j�ƼdRI?g����3���mp����Z�wZa�{Ӳ�c�>� ��m�:����b��2%�Z��S�
 k\(u&LmF.c�!^����K�҂����3.n��땻���Dz��<{H���ne�ST_,�<ע��C.Foa/G�:Xt�&5����M���È[pCj��#�8y1A�}>�@�Sθ�g@g��/��H�3�!�[�%���X���;�Qt�5�peԳ�>�U�u#r@zwoJb��˫�]�=���V��F���l
6d[�c����]oX�u��QXX_e}s_�& ��+��k�>�P��{
��Ǌ"u8A�C��z�Q��]5����a�#v�Kr� �����"ϰ`�o]������)���(:\k/�im�>�oH�bf?�s n�č$Aʋ���}�h�e�"�`Ί][����]E�+����ӭt�����o2@�z�4� .�r������ڤ��fЊ�!ڽ&��۷(�ӛ :�@[�a����*���#�b��6ܔ#Qm�6��nh�8z�V�No�LԄp3����"���jT�n��>��3���O�V�f�܄v�<B�����`�
�5�,��d��܇Wn�<����ۃR�Z��E�����fH�_�����d�ݛ�����qs�_SVN���� ���LmH����'��
\Q�3�t�.̍T��@o���\�߁G~�0/�����_�	�J���8ʘ�s�'�Y������$Tc��4,��{�,?Ʊ�eݤA�#3'�C��.�)��U���_��?z=&+�v�i=�$����V+��x��UƔy~�[����P2:.��e)=�q�K�=�-�����Q��Z�D)���n
���2�q����0+(�mv���7_�-�!&">O�Q��Ld��Ti���1�㙅D�w}b�)]A���W��J�Z^"��:�X����'v� ���2�`���f�� ��{n�R:�9j&zLy�������B�<m�����a���C��/�1�to�0�'7�n�V����+����"�EY�r�g�o�dO�.J�x��/�"�\gJ�̛�KjS�>%�0o#y��1��F�������0����S�ꀂ���)�FA��z��s�?;3cf!�Y��!�s��D_��{�E������2�l(U�(x�D�6���3����!g��f�x��y|ۜ�!�>8��4e����#�"�E�����^E�2p�Nf��_���0����_G�Q=,���F1��n���{�ݨ������p�~����Т���jd�C0.9�kp]��U�� �f���03$�T��	�ލf*q�O�k?X��H�� B~�#�U>�Z��Gd��(i�Y4�;�e�H�ge�Ð�m��ǖL�}E���2��Un��!7�f_�ˡbN,ta@+;�OF[�%�J'0 b"�:�ε���$8�������97�O������RM׬��h�T�s��)5��_�6�iڦzG�D�5�eXԳ�Ӻ�<M�S�&:���ToŎOd|f'T�I+LX�^ �mZ�̻����2Jh��0���7!���Z
��y!���3�����?�o��|���2��Rÿm��L�,ﺓ�y�u��\(�;/��5���aLp��������q5$�*�ѷ\�`aM#���OK�E���i����`ީHuu�3��Z_e�wЉ�}�)��ftu��	P8���Tz��T���'�Nz���tS�A0��9O�%H:�A$�����r�|�7����Cy��B���'���Q^�b��N�*�5.{�9�T��V�8��Q1�j��a��#@�+�vk�����Ä͸A�:�'�����G�p܁�P�A�;K��\Yz��l�.V��|��ڬ�۩;���I
ʡ�~Pc����Z&���$� #��n���1�W��e���!��Ce��?�,t7ɍT�a�yR����W~�כ���vC"b� �٨���P��do�.��>�^�Nc��;�W(�Wׇ�6ì��0q��=n"�d&4ߊy���ׄ����˚���h���7dO*'GzQ��2v&|jm���\���<6H��8�0?r�^�omG�7�=��Ap/��iV��:�?ֲۛ�/�* ŏ:�u�o,�*gJ��J�}
�*T��z�d�@ШL�O��Ȭ���
���g��4���q�E�X��4�t���s�,
s�%�똝��si�vO%��[�2�+��'���LJ���U x*-���1&�ky��^u��f[�X��/M�� Tϡ7B���?q�0�����=���]�`m	��%ޜ�*Ң�$��`�KH��CL񌛍�R���o-3�����Q벯`V�"G;�J�P�m6Z]�=-��dz�+��fqqkH���1�x�,.��q����,s��T#ȗBS���l
\���O��S���%��$sD��G�`�C}� ��o=��4��8�~5mllڍ��xR���#��+/r����EF�~͞���TI~�+�����O��1�284�۫?jN����F�ck�8���<>���Q����4t��᱕�����q�3�c�Vl�RA���HY����+�.��H3Ղ7�.�iL�h�O(K
��]��(����4�:mXG^�	�+�W�
*̱�a�]��5��_C	P�G_1��Z������wL��7E"Ogp9 R=��+nWcP�	�����l!�pXN�cɂ��Χ���+]��t���g̍r+��F�h�%�MP�_�۟o~�G�)�~o��!ɰ.�/�W��)�w���^�; [�ݷT�5Ԟ�z����6S�·=�� ��i�,��N�����]�E�$$Z)�����Xz���z$%¼���iDOot�7D�Ua�#����̮58yuJ��|j���2d��-��\įG
ت"��������B�s68}oX�ņa�p �'m��cq*+�o	��B[���Z�?'E���h�3���ۑץ�ǀ�W���]�N�$�����1�}]�>��o��ʎ��#o�c��rB�Qp���Dp2���V�I�g������Н*8��ӓ���g�=��k�v%\�����NT��
f��
,rp"�4bC�����J�i&|���s�F�R?�E��J�_��(r�3KW�Σ�:����%�\�P�݇�����_��r�_��Ʈ�9SЀ�����`�����5�R���&���{Y��y_�x��m�f� 
�"@ۅ�Kz�B�K�"�\0s2��8��7�KղHU��fEu� �:��89�-l~ܭ}v�1i��-&���}+94D���Nt"����-�tuj�W؆�<��Is��f��b��c�������|�BJo�Wt�����4��m���{�������uձ�y�Λî�I��������ӝ)�(��ԡ�<�,��U8�'�v���I�u3�����k���Kq����|
��1R|S���D2�5	HU��]YAn�������k��-���A8Ĝ{��d����S�X�y�l���'�']wO\��ԇ����E��{����h��iL�g�~N����~���)�qꤏ�>^�k���])JYC��c+f�jj��FO�o;�³�T��Q�4<��@\�!v�c�V;V���4ծ}�Z���# s۰���e(��3��&ȜM�@�e���f��I��o�����f�����2��|g-���`1azeMAQ�&��	�l��3�)A��?�0����f�N��Ǒ+7w~�@S�U"���1>���c��˷�u��D�Vw�eć������hз N������F� ?i��~ψ	�A�9�=���P��ؿ6M��H:r�X��5i�$nX���F�g���tg���d����>�#,�L�:�3��˃�LN�U�5F��?
�����Q	 |?�ej<��^XB)�<��J��S}�Z�$�ʃ�}v���pZA쓙�U�ZQr��#���W�
 D�j�'��I�B��*�	Cs�ХqN8A��7��9؀tI��i:B�<G�;C�#��=��Q�.���V/"�ywiq߷��
��q�7f�3ȼ@/#�������	�fo��$���/���g?_%;�.~[Pǁ��5	���W1X�0�L�l�V�r#�ɊD��6;ຎ8z@/��n�у�D��(=������ҹ�	�ǵ��%h���7��D���gz����|�:����5���D�2,ce�4\U1�A�qYBM ����z)D�>�����%���ދg���@��
Id����=�!&�H�l�n	�ԈjY���������Ϧ/P���cK�L	XE9@iZ����[�r���M�����̼
���=�� T��?���ڒ#Qu��~,��&�j�/$�2��T P�_��kl�},~ �ִ`�'N tmJ�Q��s6�L�b�4#�j;����l��i%{ʐD���	�~z�RL��k �4=�N�n[s/���S_��{��W�&h�T�j��B�w/��� O �`��K�0�/M�W=I���>�C~�6C�Њv�(��B��ų��~��;�y�PL�c]�dD)���`$T�艍��3B���`/V�?%b��&�>i����	:�e�ʰ�7�/�|֤P���lw*�s���#(n�2ZRX�/iʪ�;l�N���4:A� &7�ɭ��� C�A�����E��� i����K�O�����n��+	����`����T)c�k�?bPO���a?6 ��|��S�}Z��Y��2Tl�h{|�w
��_�߫�b6wRb����q�$�����$e�j�G>c<�8!��AX���b@�&"����� 
�\|�pw*P� ��E)|�^�Qp�2�ջ�E�^O�U�n	�#��ߓ��>�l�p;�ɀ`C��Ճ]O~��*�D�E��Q>u�&��#=2s�ޓ7�G`꠨N]cz��������T���E�_C^�(���R����n���c͂�V@x*��� H��`?�B��"f�l�2.p �UA-�G�%�x�����O���	]>��Le��FI�+��5D�pɤֶ)�\@�=wv.'�=y_�\M@���ë�h����ė�x��Z'<�ob~I���� #&��p��V7�Y4ZϠ�	�������::�B �o�a���, �q4��l=*�ke�E�K�?�Ǫ�s�+l�|�Ts`v��y�#%����Y؝���9��!_�)x���U�
!��yU��rL�
H�!N5:��q:���F� HU
a<K�;'��{�N{Zb�ݽA|}������(]��گI�棲2����Tg���7B=bS�\<)B&	�R�ܱ�Ž�pfک��n�֎��6T'����"�@�#�a�+r�#�'x��c7m0|�ت�&��+J���Ñ꾐��ټ�����!u���D��0��	s���b��`MLN���;��Ie��=2k�Tm-6�5^���f�W3�刉�����ӷ�y	���0�� ����گt���w�+ΛǑ���v���%��5\)�O�>�H'��D�Z�^������H���G�٦��չ�x핓�,�6���-f��)�%�o�Ƽ��6��C�ЪX�-A��H��/!�+��F 9�'TE;�0�� �������
����@7�$�1y�O��))��j:������6kܤ��C�(�	��M[����a^���}u��A�n�jM�n�䪟������G��60�B��4��AqvՏܛ�ko�� �f�������P�f]n���-�3� -�t�Ó�)<~.l���Hu�n
���+��/�[�;��VV,�)+��.��"�3�#v{E+	p-�R <[�� ���M!3��L�D�%�����q��)���t\��ϧ�3`:aEY8^x�9�ګ�{��D�z��%x�%��w�]�*=����E�f
ٍ��JU/�iX�g�|�'y��E��J�d/S*n�W�\6GP/�|����G��U�}��3<Ɋ9 ��r}�v�]��v\�9�=��rډ���cc��$��>��MX$��5!#L�;[1r�rhCODL7����x��<t�Ǯ�E�dP�����筰2�x#q5m	�`�a�|g�}�F˾��x�M2O�8�<1�
N����g(����g寿f��k�lk�4Ҫ<�ش� ��J}w`�Z�%�kul�� �#���.�t��C�k�Њ&�}&z3h����a��0of�?;���4��{1L���7���(�\����h�hC�񧇪.r�����|@4�D��i���Z�Nk��P'�lAȒ��P�2��nLM�@��k��H���c����ԝr�ٱ�G��0z����[���(�y�҃����S��\���V���:%)����Μ�?6�5�}{�I�K�9^=Ӌ�9���L�&mK'�k�Å��t}IYY�����V��=�bˬS������i�<S+�p���Z�8v �\�a~L�;g`�su��=C���d�S�C� ��.�p���Qn��������������O%qK0 \��=�����!���#h~])�8������/�-|� 5^�֙0�N��իl�Q��UF/1�#�hʠ�n6��YQTҙ��>���>�A)b�JǑ�8-�Q:T�R��o2�Q�DՊ���_+t"�X�Z��ΰ���KP|ܫ���t�kQM�Rԯ��5���L��J*�y����Z>M��^�#��$d��'��}-c8tqq��C��(NΩ_*u/y�M+P`�������b�A�%~���O�T��1��NE�%��J��aDJ���s�������)���	hO��r�QK���� I�d��<�<I��-�m�z~|�I˚E�E_�o1��6��30��um�x�~�G�Dp�<'�[
�谻k����\{�� iņ���,�ˍ���;Jm��Y�na]���]j-�%��?�	It@�4"��\�3�,Xy�2�n)���|�������%�9Tg�K��8�Ux������PQ� �R�M��άT�͈�o���aw�����m�v�ׁ�����ߖa��&֓�>9�3M�3)������[�x1��ԇ�J��ԫ�*��1�������'W�Ţ�1i���iv���n<|+������Q�n�4X�q�nG�����{���hVk{q�A���q|O{p,��ʞ}n��K�P2���]��h�aG�Z"�˗�;E!���_�|�jY���%	CÛ`�3�V*�61�����6dÑz�b=9��d B=j�������*{<�TY5� ��o?��j��=cK���7����= �ˠֺ0��mm�.]�-��]e�3y�٩3���ه&ԣ$1�0b���@=s��;I�O��U����(�m�'�X��TA��=�����/�s�	~԰���gbz@u�a�ab�(4�1�����ȩ��6AG1[�ǚ�;��N_8kz]��$:'S�)_V��s' v��K���v�l_��che�O�"N?��9�R�_�w�d㓪���z8�W���{�^�b�ͫ�6��0\ �D���nP`��tW�&�oo�J��\��?�5 �R�G��A�ɕ�o��z��'^��_��^������Ӟ,\Yg�gew�e<��F�Rb�j�,z^u�#��>�Hƾ{��^��������9��B��!��-@8��H��b-m|�,%����u�_����"ܭA��&�\8�f��nvu@S�B���
�Vt�=hS�y2���x���ʯ��e�>���>�#6�hX#���m^̱P/�IOA'���M�<��a^O���ߨS~|�}r�t��;$��sr�JQݷ��%��rbo!����F�_Ih-�Pr��n����h"�/���bZ8���;��ޫx���;_53 ����[Q�]Ef�<6�O���0�ͥ�juW��SG�"ᚸ_@��0�(����}�\�D�e�Kr��1��*��T�{a-��MǮ��� M])��v�٫IWx�*���ͫ��E�i!9oܲ/{�CqE��M�5L�B��� 3�S~M�{��n��$��p ��p^�k��,�7w����~���P�נ�����a��S���g4�S#�����B�����e�`�_����{��3L���#r�F�'<a���l��o���Ċ ��R8����Ͼ!j�Q{��5����?�6��o3F��/F��m&ʹ�D��ZA�h;� �+0.
n=�~O`D_��Y�T	�O�m��w�ݏ=}*j�De!76��״ߚ��>Q��R �j�rR���y��MIkf'��;Z�e`���cB%����I�ػ!�8xU8�KQJ���̻����&$���S2a�헌)��H����vd1-8��!~�2G�E�B���g�b-Y�����i8�[_$o��0�E��_B{C���Ȼ�H#�eX(� ~���uǬh�c.'�\�����۱؈�����}d�NZ�v�ڊ���I�/S��D�q���S�4q�.�X��yN�'�j�\��{��t6_ S����;T��PʧX�c9����Q{f�,(K.1̈Fh?wf�/�t'#y�g��~/ʜ&�4��DMe'
�B�:vq[��4�\�Sm��H�Z�E�G������w:�<��tT���,3���y1 Cz�:��#�y3~p5��[�ϰ��4���ժ���z�ؼ ��Lh��y�z�
���. r��Y�X!p�-�m�uy@pM�$3�L�j.c�E3ovu(JV��%���(��zxTc�ݳ�u���t17ss72L��EӔ&J�Ɇu�ؕ&[3�֮��w��y����${>����-��A|��Js*ݽ��U	�	ج^ǵ=�C�7;c�����)�� ��]n`��ڧ����F5�]I0>0Y��Z�Z��c�����%�Ô��8;���Zy{LC׷B.n��5�q����5���ø��Ԋ6y��q��U?�.�Ipx�l�����i�+Ϫ��a��c�6=S�c��	6�B�-�$���\�A�QYr��D6U�������r+�p����0������?v�\��~%�8U����!�K�~�e}���v��)��a� ��x�EJ4像�W�C��j��F����L�!����)@d���E�D�vO�4�+�aN�/W	���ȗq}����}آtd
�]�"�-��*����D�c�-�(��KL.��A�NF����� �2D����ʫӫ3�D|9:��'�Y#R��Q۱�G�,�.�y�/
�� U�G&;
�j<������9a����-|j�zK�q��RPױ?�9�ز �0i%z�q��9y[���6�ie�o����X���D�~�_	�K�1N?�����2����O���A�r��2a] Z�$��k�?5�+�2)�Ѯ�N+
$ژ]t�I��n��ʩ���,@�Q,Mp���S����{��E_@��jzO?��<p%uy�>���K����k�K���r���e�%4��$�'5tS�!(�Ć�4;�l���o�/��$���~�C+Ŋ?�P�,����3�A��U��B��:�1;`����,o��"ލ:%le!�@��ckY���!$�!ԘA��������x�)^�� �ҍ�f��E��YD��.z��u6�K�K�/����A6%�0h T���䳷	��ݺ�q��
�djnjC���=��/�mp��i�PڀX�-���P��P��w�%�LC=���\���b_\U�K֙�J�F.�)�G��;��fM�t�>�vS<���k��f�]���5��4v�uׯ�؆�P�����?�5?��ߔ��&f4�굌�$g���D	q�4.�m�b� �����C%9�5��lq���q�w�?����}����3kM�8��+o�tK-�T�^{Û�p��;k��P�_�X���^��$��6od�Y.R������W��O�o��p8R�?>��"�_|1��DxC�@vO���Յj���I���3���(C6X@��5����τ�5���j�8��Y*�7�_�>^�"ϝ��E����*����4��߁�<'�7Pr��Fz5�	�f�:�6g�LEe<?
�,����1���i�ee�;�6�_�`;�M>;��]7O4'>����H���>3���M�i]��g4ǭX��pQs�=�|t0�������<ܕ�A��wɳ5����[Y���,�����L*�^��w�0'�6���h++� W�4-+�pu�=`�ԋ�s�U'��d�{� 	����ٞ����Zt�����w�P}('\�Lr�[�*j���>P�ڢ�$�F�P�ν���޳ Ł+ ��QE���rS�n�ڽ�S.TAD3�E\�/� �NG�%�i(������{~�:��=�	᯿��)I9� t&G�w�Fi��h$S�z�mჲ���1�N�'�F���7�Bn���3�
g�5(�Sr�i��a?��84�
�a��!/"�W�O�i�l��l��E�(�.4���.�%�\|�����ى�_5vYq>Ƴ�H��@w�-�p�-�wD%Uq̨���X��}'<�F����y�;Ի�yߏC��^��Wb���@q�J�$�C.H�O���B���P�|��l�jǣa�K�{h@��|�j����7�8�.LKg��!Be�O��1�
?�5g��zS�@����;���v6���y��t˦�ڻ
�����`@+a�Y/����.���[Ӯ+���X(X��n���"o�������
�=���{]��G6�tD�~�p��S������rŲ��
�[FFXi�k�BPyd�0��se�	���j�Yrc���-k�o#�*�!P}jɦn�{�����!��%��>�|���?�TD)6�>�A��|}7�GA!t��>0D��
P����j�)-ܙ�X�%|<��7^���VJ*�k�u��Z|[�&�ḊmvDٝ�+�aKbGr��^kX5��s	����6($)�g��$�-�^�Ňe;(�Čn;#h(���ԅ}��􊺽�xY��	N:��nJ���;��y����uD�qk� o����-�GO�ݳ� Z���SN+mr���}*;�*�E� e����h0���^�T�G-�ڂAv�!��Wk"��B�N��u�uA�m�j>1V�v^�q���1��`m;fڃ7KZ�Ҕ\y|0�4�6˧��CS;:U�H���8;]�������P(�H�V��z�e05���?Y?G���#���"��wRɀ02��9b�_�]2��=bَ�(h�H&��5'�J���;A�fJ�Z��ܑp�z�����zuq�g���z$�Қ�	�c����"e�,��,|�I{�aI�w�"?Z�S�/̅}%���Pr NY��^�Ռ6Q�O�`��
�2H���֫E�Gu��h�ԧ��W����}֡nP���b*|~cot>���9>)T�1������)�B)s}�?+�kY��}����C�Ɨ�mN�0�=|���K������?H�Y���L2)*jD�}�~�ⅷ೼������THC�S���S'RY+�Rϯ~́���q�p�5jo#��aB@���@�$����s�Qf�O#���a�sB ��ݸWJ�8<:�5�{K]ڔ��A��2��aV2��Gm��c~Ђ�6���j�/�I�]�g"�o�S����	�'��?LrԑZ���D(����V�?�~[���iJt�k�n�ehVy����Tb��,Pv��Vc�Z���
1�&K���%K۝MH�{>�w矾y���y���a�U�PK�»�dX�?�t���մ����7  �p��x`^\ZU�����j(����hFu�ND�[v7>n�{��6K��9��y����%i�>Fz^�38 �ZY)�����z�DV�l^2jμ?|�q����
�o[ol��d��ϒ@O�Z$E� �7��A#�j�+_�Ns�ON��u%���V��߹n��]� V��WE���\�i˼ș�}s�Ax����c��mo�%o\v$MA{ ������I�ƚP��a�X�;�5�8e��,r��7�E����	7�Q�s6�� ������h���,���B�aM>He�X;_���L�Eip�85a��>�{������λ�'3�77O���@��M��w��	�o4��j穊N��A�W|�TN��*$��gٴf��[��h���C�}����'�&1�8�ں�ܘ��;�8A}������\j������9��v���U�?�׾��I4�o���+��_P	WȇUlܥ��~ӝ���ʀs��?�|4>6!]�|Z�Iο�)m�L�C^|��Yg�(��P�Ho_3_VN�K2K�MMx�~�(Wy�w?���@`L3M5QɡG�Ak�N\��a�@k��Q��E�4���9�/qq _���9H]r�7�N:�6�D���"�L4M*���׎�d1����!`֏՚��MMĜǔ	�[IsI��&�C�2�?&�"�̒�ԟ0׾�¸���Y�2�y����{Q.��7U�{$�A��� ��"�B��Kh_��p����@���"�Qh]{1���[�$X^�
(R�2yS�aNT��Y7 �]ӝ�Mb���O��%�8+\4����T��8+A�g�y�b���1v?�M��;�}�ü����x���ZR�%;E9 uP�?O��G��^���	�qH�B}Մ
�3�S)̳�+z9�2���qW*p�P�d�+*�nr���.~��B�=Ώ�Y��<��O�Ǻvg|�7�ƼQZ���+�����s �^�=1l2���mm�6�$�ӏJ���yki���yq��2����_���K�2,�ǰf�m��W�dp٬5® ��-��0P�K���Y"@3k������l�y�9�g�W0袝᷎��D���UV
{�@���{��MEӏ��QOqm�
�ЊE�>xq5�st4)�./�$Il*3m<V��(}H��Y���cٜ6��M�@J��m��F��'���N����ޮb{*�?��`�6�=ե���4��K.��RXG�����*I��iA!	��>/�*vW8�Iߔ�rS�:���xFYoM=V|�^�;��9�ކ�Uf`���h` g�՞�F> i��Z˓oj��q��Ϛ�������wkg/���M&��m���nRj��;|�Ju��E~ΠQE���X+u����uol?�ׇBm
�_� i[S�;)�%�媅K�E����8'����ȑ���G�;��٥�󎹺�ܐ���2"��D��|MJ�L��@�#>��Op�% �VcV�Y�Gn���`�E^lR���"RW����̰1�T}��c���sI�|�Rh�.�ө�}�ߚM�`E+�i�{�[�/���G_k~p�I�fN̥F�c�=vT4�9u���b�%��2 4W����~�0@��yـOHl�s�9�c��Wl=��<��)�wZ��_��
�Ұ+c�g���3�Y#O%���%�?`Jl��V,�:|�v2Y�Z�ܿ��r=w�_�?�<X�®&���"I>��mID kb �"#!���Q��A��T�ߊ\�s��QVK��~�_�]{��@
�>h����C�hE�G��w�ذ�p.�Sqm6��1�@��e[VS�!��Q�DF��y�o��U�חҍq�A��"�ad��j��r��4�bL�8J��� �e�~V� ����\.�-9ӧ�B��R���xv_���>/]֡0���Ͽ
��Q�4�h�#�k�|�V�[ ͇��ȟ�$ȃ՜�����,͒��=��ā=�N��0��W=�i9$��3��y'&$��rn���
�!�Xvmu��o�ɺ��5\{Q�t�	���,m`��!��"�gs<	#�H��J���n	�D].{8�
_
Ƨ{�eAgH�����/�ζG�I9���6�i�-O�E��ˠ�����Q���~��ed*s��C�\|l�x�a��~�U���ߖ(2!�I�x�٪�N��`q�T˿����+o#�f�!���K�oT@��F]"�\Mgvsx��&[#E�?��^�LBg:�[�:������A��I�8�O%��o&�� ����!F>�Xe����~��ҭP�O໬��,7<�u�
|�]����т�:��`�M��ڄ:�o&~`sd,YyB��d�Ju[qE���-����c�������rR����	��r,�>Lc�>e���OF9Xy��h�b�����Rs7:9%��K�}��yL���A������� ~�`����F}�kW�J%C�EQ��|E�n@w��5A̕�p�A)t������t���������6y�K�?!�M* N�MM|?��7�Я?����)e����L���[&���P\�u�r[�c'�^�o�� �6�gi��$�WO�_��
��!����i���deK���EYr��M�%(�a���U�<0�q���6e�K Y�/�Ok��U�8Nr�hw$�+��<��؟���5Wϵ�A,������ �����NG�<����.䊶2�P��E^����В�d��i$�Bi�j���\�:�, UuzNp�󿡶2��q�R���yTsv��h�8oy?�u	�������a�d	*e�Z%ˉC�9�h$�͉���/���>��s�eQ��l���� a���P�^�+�8vN���"�W��BZ��x�n��jmζ��x&W���1M,_�	B��2��+���'��~�~ā����R,<�vl o�x�zy�_��1�e�M��{��rHmha�I";",uS�:�{��y�s#~h��H����Թ�a<�����FoĎ���!duMG�!�hj��L�]_nG�@e���$����ɛ���,�8Σ!5 ��G�{�{G]H�w�N�$^�����o�\�j���;���=뚨�S���+q��o��Y��:�
��! Ԭ�����IHǜD�f���g�$}�Rg��
{O��I)����ƀ�*���\cQ㋰�A�o��p���3'V��h�1i��*ܿ��$΂����n��z_fN�O>-�s=��#���8��1��o���}�>&aU}��.���D��@a�_ۡ�E� �*�i���(�K�3��^��

D��2@dr}�Őg4~K��^�}=�i��#5��4:��Zc����\}�]��F�����,�f�`����M�B��]�'\"���2�|t�@��p߇�(����/ !5�SѠ�&i���sƼ^&晏�9�O����֟�Xf�2�mY�m��u�\x!�Xsx��ތ���O�5��h��@2��#WH��0کT;�{�~�����Zu��_�8m�93��S�9�%����eF��ڹW�'5��9����R<Nl��j��fA]�A�ys���_1L�6��4���M��'��yEC�v�`���E1���7�:�E.�_�O�����Q��6`�S,�NF`���������l��nd�p1)v�L#z2���.�~��AB�Ϧ�~�u�j�2�-IU�鳖Y�����o;��r%obE�{�I'�R}�]ݝR!i\�H������ה��o��e��i�?������[�m���}1ӗ��Ev�u<p_J;���z���%c�EݼXU�����(�"��vվ�+h! ��Zͮ�)8Y.Oޫ5��^@���SaZ��9��{�x������R�Kj	T���y��O��9�����.�BT��7t\������w�&��{s�Etޗԅ%H���\tDc�Tp7!0z�ga�$>v@oJ�\
�9��δ�31eQ�=Eě���F�!2-p�~o�J��m�hu�d�*$�����z�M�3�ǟ�O0��]���&ܓ^���ctC-||_���c��X��Lg��Ve�>�M�\ͯ-�=�{��F����ª�ܓ'�m��R���'G�����3w��WL%кU����_S)���������J���2���:��o�b�Q4��b�4x4�1�]E�|ll���6툞��]�뵅$#�q��Uk_h�P܎h�dw݆����X��~��5��r���w ,U�U׎��㞕/�[w."��R�{�x�T��_�Y�O.�5�L��}�쮚*�AsC1l�Zv�MrĠ�{e}���*��8�_�G�.��u���\��4�3goN����/�$��a
"���P����c�7��C��̠��f�\6�/&�H�;�ﵧ_�|ؤq-��k�e!�E����5�N��8 Zd׊ԑ��B�#�4Q�'j�l;��`)D5y�8<R�q5�R�5@��Ϗ��^#�a"�M�5�φS0�"�_��]�:9P�빑.���1:D"���|w;�c�<-y��n�1�"��B�pIA#9����B�X�d><VJn����r�����,r�zk�
��}���#�b����{��ciZu��NEw_ �R.�P5�&��O�0�d�ʹ[c��^��� �\fխ%�r�d	��� ��,�li���C�b���Q�ОQk���r3D�ᅜ��N�
���{x����Ju�oR%x��´�����ga.5��q�27�u}�������:b]� �dx�b�&��{ư��Hz9��y�wk�o�^_yMr�dg��e��D3��&t�:`�1Jg<��1�2@V�8�t��0��}t^J{5mźR ��8?�M���B�/��s߽G�A�ƅ��}���l�p�'?b���&:5�r/��Ne�����vB�?d1���x�X\}ҭ��:��z���N@�������g/�4��G�y���0�� t*aݥ��^[h��=�E�<�]���3/��ؤN{�Z��JɃ r�59㲗"��^H�;��9;�.�J�q&����]H@W}�De������T�>r'�Q� �}�� ev5�:1Fa �[�_��O�N�y�R��Y&�n�<�w���S�"�e>/���9�bo���3܋����i��Dy���Y�0XL�gF��!��0�Űbf��"�fk�n��(c0�k��c_q��TMĔV�|,HN{$�-����(�i�Ԍ���i��8L�y�s�`e�!���Ք��Lr!v]���@�1��A���7���1�+68���|���u�	�����ZT�a*�[umTm�%���Nx!3KN$����ɢ������k/TY��icuF)?wH[E�n��@8Ki� �o�ni�ų��@��.t�0��gQb�5�h����HB>]DBH�+��U���gH����4�x,A�$p+kMm�OP^��e�`]��]����G�ա��N�J�w2�^?r�Oq��ё`�Qit�;�T�^�N����cB]�Tx�.ls�4p�4���S���;5�*ca�on��� ��r��"L��5�v���{��a�._�&t4(���_]��Zxu$�DT�����R�J�t\Ն����4��(��G�QtY@�B8�G��kV#��ի'���:T�s�ē����G��%o��M-�]1����\$O��7'D? ��u\ ���E������g��"|5~�Ch���������cj:����3�-w�^O���%|��}���#<�VS�����Ad����{ã�	R���%�0�R0�C�K|��bmtc����mL9�`X̆�n�G�+��j�e��
��BKu�[��a�1����Ѕ����ML�{R��S�� ����"�ïʚ��_F�5��E-}
R�.67�N1�,}���H���_ٴ53(��N�V!�=�Z��f]�ΒC���+�?��u�B�lZ�W?|Z!�,�~�疽+�ד�[�V,�����r!"h����1�ˉ{�~.-��Se���ƟunR����w3�H��||a����z��F�G	����܅�]��)�D�̳��nN?�PVn���j����@r������w��V[MDg|������p�?�5LJ��1�JKKm|N�#} 
/D��0JS�j�7��`S��Id�����v!0_./���{��D��+D��~��,���7-��j)��mk9��¶��9����ߔ(�9D�ٛ�E/2A��{�Giw�|���<XC���ᐟ�A;ِN^g�=<�>����˽�/�EsX%�O`@R:��*�h�0fcTh�P7W���G���m͉�U��d�l.ET����j�u�ҥT�`W�m.���-����j#�f�X���nu��]M%���!%>Y�'j:�B6a��Z� �v�	�Z�ҿY��3U
�@�j�����w�������-�sr�m����	��f�b�*�h�@ŗ$3>mu�,��祕����?��J?qr�r$Q��'w^�=�E��=�Z��v��Fi)��ٰ�d^G�^ӻp{���ՙ����e�}��j,��D6��؞��! ���
�Υ�&�O'/�4���S�3�5���7ꁡ����0���:��m5���QJf��LR�����}vq%:l�xp�a7���u'��78R�r5�d ��f㧼%`W��n�7p�|!�ҭf*/��C�oܖ��9���(Z���D�(��_9�=/AS�����U��ċlk���L��uF��iu�j�K�/�
�U<:�5j�5
�H>"�bE�ē���M����#���
���<�r�S6��׏�[]�v6�G���?\����6��E��Ty_�G��x�̓�۳�~���Q��u<�Q�?��S�-Szd�?���Cg��R;��6,��7�|�-�^Z�5�Sg�]+ɏ����E7�I�g��C~��A����Xz%�<�X�k��	����@y����j��`�8�ˆ��◇���k>�^m���{���� �Ro(c��~�\�p�rj I8"EG����|C_���ȯA�@U]ɱd���Iɴޛ��"��V9����U�Uq_�m����=���ı	��L�՝9�eO����,�6�8��*��0��b3��"h�G��$�;"�uLP}���ɗ�Y�"aQlOzýC �2�6��\1P�\,+OE֜���L�&���]Z���7|z�"�¯��s^��u}(�DD�Y[?^U�;,R�8��k��kZ�x*�w�U���kA�r��������_@w���f�'�6'�^�	Y���˱����J�
?H�p����Z�I���0���&���mD:2m��Ów�Vv�)"��q[�'�Ā�]���̣u�O������|��j�:�V�!E�FضM�-C~�� �J.�
��&ӣ&�ZxBa�%X� k�ɐ	RfJ�F�&ց���t)>����1i��y��Hu�����A����H�{�D��t�t�bf��y4�UW��*�Ut�f;�G��̓��M�H3���b���"����rSk���t��ţjQ�F{rL����k�KU�2��
=dB�0�%�
���\?��T!|"L��+���ʠ�	��f�W�2v�~9{�C2��@QO��H��Q���rs�/�jߏʜ[��Va��O�D�\K#�榺���� ��4F>r�C?��u�J~@��;^�ي߶Q"��CKE�NU���e@���Yu�v)%�1��d��C�pZ�&��>�ֶ́)j�0o	}�y��|Y��pU���3`?��\���t{�p�@y�,tw�9����M��ھr~C:�8 Hߩ�@h4�B�����k��ψ�ߎ "�=�� Q�)�6�ard[���X��Y��%%]�(�jWs�0��Iw�5���Q�C���͖�P���d�8����Rc2uK-�/SJU�\K�3�KݘX��cNKLl={.sH�3E�n�
�`���5�y�^�����)
����J�{�	�i�a`�<�Fv��jFB�q���'�ׁre�Z�p��)8�N�����{��X��3,;��#>�#��ю��3�}C��_,��?S��`zp��V�&�k ���?k��4Z���x�1�u$u�?�t����m������g�.�D��J��Re4�&���ѹ<5�B����ϭ������2�U�����B*�cY�o�ژSƴ��g������NYt#�PtjF�l�G��u���,��-"���Mi]�]�h�HJW�yy�O��8�FW����qs[�v�fE�g�>�\�����?��^�R�5�}�b��Ka����|��zp��b������SK�9��c+.��W�'ԝ]��m,��
����U�ѳ�Ͽ=o�	�V���Ȥ�N�f)��db�T�,��d��J_�U�s�M�Jb�����-lV=Ӫ	�_��nՒ��rĔ��L�u�yǤ��d�E�
B �*�@Ra:��;2�#��F4Uk@剮:�[�#�t{�az$�D��8��=�gD���.Rq�r<�R"��i:�����P�[��:��n���Y�,ի=Md*v|G���;�b�K��ߔJН�����_��Ee��pP8�6����DT�z�c�9t�R�@=��Ƭ�]~A����8h��.�owo!�ٌ:�K�'��,���6�vM���H呟�U����Z�ta��LF��g�+Dȶ.2��^���� ��͂Tg�Z��
9�"XM�Rt�4��;f�`�϶&G�Ċ��7���!E=�9,��4噬̔��Ň�E�L�-wg��P�~��[9�-.�[c���"���s,8�sbo<�7�J	.���R�g�b[�<�/ƿ1� ��{�G�h��&���� ����8�
7�3�[pہ�ujGȋUX�1��Rm�&]����C!(~��}��|�h�"'�H����f�?�8�H�#�@�۱��"A��˃ <ٛV���kA
Nh՗����� � ��0Yʀ7�jT����VpP�J{ `AX�������u.�q'b�x�s��YFξOa��l�HbA�����Yw55Oǫ�1Z�b��L��dk�8��}r�?��k���A���L��P��Ռ`��]���Qq�%r�ur-Q�\��T,I��"�Z� ��c�vu��Əe�!bپm��I�B����r�1�m�_$��1K:]�ᘸ.At�{ ��� � 8q����_�����+AX��=?R�N����ьH�U���~�zH�ώ$P�[�^Iӽ��/��ai)���G��W�i�/��L�p���������@S���N���Ҫȹv�,�Ts�Y�XQ)�p��:�S��4���;J������j��8�V1'!4L�7�>Z;x��-�HF�4���c�僷OH�9�n����wɫ� v�/��n�l�]J�9�=�]ѧ�~aV�?�}���&Y�+S��o�FZ��҆�ST<�2�;RM��l��H�r�@�zE~iM���|Ө}_WB�-�Wbԕ�6+3�pZ�|B/Ҧ���*�����j'&-�u׮��hqVC���ז�˴t���P�T��.�Sh��G���Ƽ�Ė�����=������_C.RY�J�,�D�&�B�i�cY�Њ�=v�;[Lƴ���6�P8!SPg�XgںM�6E�j喣f��}��=0ߝHc�f��O2BG�g���qe��-uk�G��X.�I�kDi'� Z��(�1��tB�8�	Qam�7��w���%��9.H�����K\�~Lx.g4!�LL����W�r��h�ש�z����;V���fh�WTx�5^��.��u�x��w6%�v�u'��0�=����q��9� ��")�b�N����a�el�����B!�D�zd=W2�����t�F)p֪�~S�{P=�H2��>�m'�K��ϝ�/���D�ȩSE���Z��V�$�e���ov�W��זr�����mrY��}i�t��{�䳁��n}_� �%���ik�vN�9�~gkE�֭L�7+��v�u �[����k���u�3W�#�'Z/ݛ�H���x[zK��&2��m���QY������b�v���&+q��]!7��H|@�};H����<C�O�(��(MWu"�}��?˿��Z����J��h��*��>ԗn����Xsե���\���y2xLNǌ����Ya�<{d��i S*�Iǒ?E���|��R˚�][ e���_��?��텍iQ����VH2F �X�Nֿ'<p��PX�� �e鲗dr��*Q%�� ���y���#�;<R/QK	�D�,�k�6D��Jylf;9��kp%"��Țb�*)DQ e�=�AwW�^N=�*��NͶbD�_�/9)AJ��<q���<��ø|���8(��Uib@�L$��Ŧa�-Z�P��B[_`��3�@,V�CUT[e��_�t.ie���������'�KE�we���\{V0�%P�b'�KΚ������t����!�/Dޒ��O����ǥ	/�C��$�2�s{E"s�5H����^�I��'�;��#�g�O�l�tZ	H.T���6sYp�. �{��0]CҮ4w/�CG7$����0�NJ�a8/��j]���R����y�H)+?ɮ`�'DܧJ���͞7_P+�c�\��	F9�H��2���`�Ϙ��D��߿�po��$�?l��-n������m�`jY�ҏ�%h�-?l
;ݪU=��$<L=h�އ���U�ɩ>	M���ĎC�3j^�Y�V�UE���[�Lu�&F��rH��� ��=��/�1{�<�.�9 b+e�6��_o'����G��]H�xap�$��z�9`I�R57\����vk䬓i�	A�|���8/���Ch�@JP�]>�&�7�Ĉ�1q��q ���d�m��S_�/6J8mt�^s�\fھ༖V��Re�g���{ �8~v�щ�ı�0��来hd9�ʥ��5��9Eh/���j�|о�.6�#�@�ӡ� 8��n��}�!�����o�(�w��ݕ9���@2����ѭ>kqN��R��v�U�P7U�"̨	{�`󗄏���}��(r�_�4�J�%ۀw���%�5�hD�`�5n��i���I����k0nX!d)�&
A5P�5�O�l63����|GNy���Y��5`:�v�;����9o� ȟ��+���-��jם���y*_�b�C2=���-i���
P�=߲n6+g�F[?���?6�����̡Vz��L�p�qz�-��uǨϢ����Z�g~2�ׯ'�u�n����<\�	킃{z�8pC�A!OK�n�y0A�=ۤh����iwhS�6���$�1~��h��@�aP��#�����Y	�ePmD~�[���W#���A�K��Hub7o�ӫ�A|���vD����b�越'm�*3��=�̩2�m�������Y��u�f�#�sm�x�"�XR����`���:�"El4v�R	�:� �����R�����]?cg�>Ue,��gU��c�#����Y�S3w�u�{��+*u%��s���5�^�6�1�Q����7,~~=M�����Xy��$��J��K�&��)E����$���:ы�t�Ն�����uJ�'0RJ�,�i�Z�y����D9l��yM���>N�ظt&������{��:���Lo5�sQ� �Qz��z�ɼ��D��6&Y�LaSe����e2[�� �Z��S��.��%y_�f���U�K��� ����H�R����o��<���6fQ�+�q}Эu�P��K�lh�f{\~�#�1��Y/�J%!����n�4���n�e�	���,tӡ�1�V[��ԩMHw��9��o#�N�Sg伏l�[$<�F��x�×E���Rnx\��3Ŀ-�$~,�1�go�t��V�? �cc1@�r�����=�B�En�F/��HC�z��w=M�\��&޼�e�d��v�I�s0��J�6�J�F�5�59�?7�!�ǩԏ�
��sb�\لM����s�k���Ũ�i铓0�o��L�R�I�IR�A�8�D`��A�d�,�2)��_�~a���N�K����7O�@y~��Ŭ)Y=��=i��L���Շ�k��e,��4f�Tu}kƹF|�ި��=�mVN�Ƕ6�|�'>Y�y�`�(�f�AxQ��k��cʀ�K�g�'�w�����0#�z���6~�VQׁ�3�<�\\o�(m�؏�Ե,=:���aT���n��7�0�FD�[G�@��H�b�;�J�-w�O�e��.��.���%D��9]~�Ѥs���bn�D�E�
|�}�%�C'��Ͱ�o��7��C	�����3�M̻e�������3A�$�j+p�[�c����No��)[#����UV����������:q\{�-N��.i,/]�,
S�P{��,����~d�Z�1�(��ʍew�O&~َ�l�?pQ:�MAM�܈���I���U��~��>h�lj�� J�G5f*��}l	�u
�v��W
��{����{#���iW6+dr�Q!��ʬk���5*�8�hlQ��߳A-lR�r�
YW�V<�~~h�h���7�?�V�T8S���i~�A�&�ID�K�,b��>���mGf�uo�謗T�,g�Mmy��Å=T���k\�Qh��[��9�'�9 �%��o+g�P�g$�#Мϥ����С�Z��^�Q	g��uwr���Au�R�kj4�cf��Pxس�'L��"}�p���B�Y���!b�l���a��ν��.����"�3�Ʋ�k�|, ��-4�j9T����X��%��� �yRF�@H
ۋ��*8�"a�T�>'��l�`M�Vd僶YMc�q�Yz�,�b�Z��č-?��wRײUv�GgJ��Ȯd����%����8���rZ�`�E�"�;�G9�:����&�!�'�u
flC�ДD�5��G���gaN�s�ǄG��{!�u9a����:���IZ2���`*u��^^s� ����H|tn��5J7@�Ɠp��� �gɃ˥�[�TL^��*�
�^Y�?�W����v`J�6]�2�.%�΁ҿ��ӟ�%�;Y��-�[-vɋ�o�Wr�HW'���
�}��3�m&�mGQ���{�	��@0���NEx�__��d����L1���xdQ���DS=>�q�Y�,9���J��.�������K��|@@��z�q(��#�?Y7���)ﰈK���Œ>�:7`ǥ��E��NR��(�Vqt�d)e;�Ak��iD%�2��
��oX�Y�n�16� �TL<�'�c�����I�f#��zfp��g=��&J괸�E��VTu��~�b�+�E\�傷��6-�3�O�X��;o�L�'�B`�TW��%C#83wu��<i~8`�S���f`:�7gŷ�?㫋`A�U^[��UK.(�j���q���d��O�@�_�H�u7�MdȼC:��Z�FW�˞�VVGٴ����϶"cƒ��]is���N�[�+�T��	���X:��ZN\P0U��
��,TC�C�!4�q\��zE$�:*�����\�$ ����.7����!���/e���E�:N��m\?�{�drk��^��;`�ni�$ǖ�FH��&6��q1�q6arl;�io��_�}����}������c=4�28�T��P�Mz;F�a�� L`��3�!��	��ZT��#�m�N��m�^����u>���[�G�I����H��՞�|(�!��0/b0_J�m4�ÛC2�����*���G�U�o䴴ԋ9����2��k��b��*).�׍��&~�� �_<J�TJ��E���L���nh�d"b=���q�
؍l!B���ǨG����v�#6(^�K�K_�v��1:B����OŤ���6J���O\�풜�*��_l�%�fv?��@����Wi.�7ۑ����
�*�s �c�wc�o��7�W��~h��H�[���8�텋������#���9ų�L A>��B4��kZ�P�����moa����C<o0�8�I���W\�+?l@�VXm�V���òE��`�!^�#��������%Y���Ɇ_R�<�g��V犵t�E��ĺ��/����@����Q���기
b��p6���~�b��ǽ��X�E3����M�i>���F�7x�=���jj�2������;4�S�3���.B�C�V��r�siNh���at&<�CC0����x�����}?y��"L��b=��GR��\�M�c�tF�P�N��|a�_`���o{^+Xka��е����1ăkP!];��4e�gꀯ�g�D^�^���@�J�ʖN5*}�!hi�ih �܆)��E���E�������{��>L<����!Q�[�u�����ř�"���Q�0��|�@$EWR�����@n���(��ed�0��'_e�^v�c��w=౞mp� ��[P�]6��5�̈�A�ż��n�	%��-a^�����DŮ��L���rv�f��D��j�Ic�
+o7�$G�ɻt��ݡް�>$�9�� �G��l;�4=��Ye�H�'���2G�O��;�;��~3���%s6|j����ƴ�Z����]b�~D���ە\ط�ʽ?l���hX���o2�S�f{��w���7t	�pC0��>�N��3�IU��z֔I��cG�EX=a�����r0�c< �;N�,0?�m�FV���0�@����V5�����G�j%��{��7/��Gg���kQ����;V���Fq��>Y�!��E�!! ��=1	|c*�/e!(�Ꮁ���5%~W��$ʝ�F������\��)V�!���w�+��`mZ�[aM��	�y�[���V�}�Ɠ���1�~�w�oo�#}��⩴�5-������47J����ם�T3�U^�Z ҃V�l����>b�����t&�Ơ�hJ�ql�@֎S�,�wk�x=u�4W~�l�G�vH�}����2� �}���V�"������j+zz=�)<�/lk9��`����2�47�U��+�)i��-��	x[_��t8q�h��jM��&���Glى����*��F����P3'��<��V/�����f�-8*]N��ɗ�X*��>�x��;�O��i�D��^*��ڬ�����W�Nt0 g��y��:ޯQ��/k��B�}3���}�����ͣ{���f{r�V��O<0)<���z1&[8�P�{�Uk���IJ�n�s��Hj\�m�e"���#��x�]�H�.�^���Y�B)^N� ���ex��ȱ#�vg���&#P��+�~D�Le5o��)���E6�tU[k|�"�E/o2�bh0�xiT��Y�iF�yw�Jb�mӅ��`��xA��uPK�Mhέ�����eU%',X�0�Ձ�ɽ��I�"�����;dO׫4�=?��\GlK]&��G��P�=��8&����_����c��ia�O�j���n�2f��X?�\SEskV^jlp��U�E�D�t.u�6����zڤ?B�]?.#ԣñ�I�q	�R�DB�dvz� <�-Utb�,\O��.S�M���;m$�G���`V�ظV��+7kc��� ��aJ�[o��)
7�~� sOw*�p6����� ��I���h��-�)DN"+\]�0*��G�t)��WNP�
��j�dH��]���|�Md�,ʇ6VPV�lս�T��7=)��� �B4��3š}m�A�M�hd�R֥p�&%�{��Ԃ���%����'��9]���q5���� h�123M<*R&�9hE?��]Vw4��}�k�5�1����:Z⯱�n�Hs;��z z��`��x}|�dl�9 ����<�RL%;�;ʾW���y��`8e?I��2�3PQ��:�����p5�h�o�#������^9)G��G�d�k�j���_��I�#��$��U<��᠋L�d��q�>�Ai��(j8��Fd+$��LJ�i�� ���_��0?�1�_:Ս];ahHH+%5�M��!�)VD��F��U�{����6��G�>��faTK�����Ŷ�ڊ?HK�ޓ�� a���l���u�D���4�H>����	ڃu.�#��n�S�N�F���riyt[��c<��s(��q/�:$4�?�X]NUc:�q�\ ~�M��&�5{?�a�v�y<I,�B�WA�C�F�����ͫ�W�Y�g�G<,�b����s�r�~�����Ҷh��}w�0v}��=d��z�2eߒ9\am�ז��P�K��:>���uC�5M"<��5��r<X�wf��
W��y���)�1T��WA��}l�EȷÖ�v
�n����)7��k_���c{BPG���#��0̾�O^��/BM=�@˯a��:r4KS�9�W�}�S��牑M�-ll*T����&ݢ��P=��rF��П��=7q��Jl�i���� 2?���}+�X�ٛ���!/��C9����Ó�
l&��`�N���Z�d��V�|8�|h��R!��@���+�7�i����W'��u�Z����`�R5�p�y���k��l~C��Z�(:$��q��JҨ�K���Mb���ij��曂b~�W�X�P�G^V�b��N��7�!��m�欅�<��a��6O{����║��ȋ�z/�-h4�X㳰���Ku���T�`^�Xa��CW�2c���~ό��ĺVF��,�i�����ׯ��lr��g2jV#@ꋻ�P;W��c���<tA��h#1�}.��1�h��c3;�=����r���'��uB�9�4d1Q��# 9�7�]���
�}r:�7B׃d�� ��f�H�wJ�{����D�����K�'�	�/�����|=�eQ�bJh�)���c����ަ�y-�19yվ�r�(�ё*T�wNhɳƺ�0����@?��AQ�������e�=0�O�g���.,or��'(�u�-��hk���N�Z����?<�rS)"�����f�����@�ї\���قܼT�5��,�S�\]�4�3E����}�5п[���4�g��P}fw�ry�!q�̓]+���fL�j�����F�p���t��@�w�c�'�m��^W^^�p��;y��&Lz%������%ڔ7�|Tbh	*��U�&R>����^����W�\F7`�}��%V!�7@{�8Ӵ|W��}��it��{�3���-,]�����0/�{?�T��I�,MUw�eo[M�y$���"�>���qޡwT����K>Մ�{�N${Y������S�U��k�@A�o��4J��~��62���*2����YVqƏ�]��k��R��	fp�����T+-��hQ�:����ѹ� ��6�PX��H��p����7��x5z����9A8u-8TA�
�W��@��.��#�-h�@�ޱ�̔g�Ͼv�H��iq�7�R՝���}R>̧/��8����U��� ߔ���&F��S��&a
���|aٙ�������6�IB�Z���z�0�y#s���y$B���������v���h��<�G���ΰk��<w�v�'�� 
�U�毃�J��ܹ���Y����B��(���w�3s*~�T��k�cZ:�0via��xG=�˧��ɢ��[�h�����y;�U��LUG��o V�����r�z�U(�Ӟ5���,�/�"��r���#Vm��h
�i�6;�-$;i�ׯ� rV˲q��.B�����+w7�>(�xQ�DC0��p��|�Y�I��"B������B���]f�H�\5I+���l���lW}zh�E5�t#q�2�ێ4�1,���-�R�'�ل(��T���]�=5o�s���P�A��^�T���d��P� Q;���ө��4��Ȳ& Wo�!hԞ�ya|��sb��V�	��C4Aɶk��M�Uz��/Ȝ�Xg���7!x`0 ]X��Y��Jf����� $���a�ay\_%�Hb�ю5�dc�4�8DFc1
��mG��|п��h.؎��2��Af�N���L��e���'�t�Dc]qxK)�$!���(�̷�~b�΍��1�o��8�_�B 0um�>��Q�෿{�y
����4J�~[�ۉ!�ud>��
n�Q����DԹ�$1�t iCm�#5�I'��̈́�6����>ݵR��q`x]~��(j���T�PƮ^u������ND�i����_�D�&�c�~����M�C7�F�I���V�d��]~�+�Mۜj��;TAdњ��W�^{�.�h��~�ͮ(��%T�x	�q)�R�>��4rԽY\�pY��:T�p��j:G���hA�X��g$��6���3�J!�������/�\�Y����挔�;���mz��P�aŢ+�|�{�d���N��Oj�he��
t�1��=�hx!�:.�jñJ�ӣ���.Y[¼�ـ"�Glj�t����Q�����g��:��Z�@c�$8�z��;�3[Jq u���*�q\ɾӫ�a�L�B1H��Pt�?S��)
����.�o������nh��
��	`�G6w����f��z�i4]�vR� �+R���Yj��O@+JԆ�,6�l>��֗��G�ʶ��E��Ե���FN�YK���^N��%&�ݛ5iw-���2�.�`a�|�&=&wT�%���"x]��3�0/ ��$�))�:i�Z���jR�m� �[)fQdOU�ߕ�dgr����ˀ`�[Ы-�u겈�1>��g𿍥�9Y�2*ϋkb}s����-����|�c�1߻���	�!.��T?��ʣ@��������4��%ѵ�
�ƺ ����C����R/	%Aj�1Fĥ��5�g�=Biqb�9$V���/�ϡ���ح�j�IF��Z���a"n��sa'm8��?e�S��ϝ�jZ0��b1oã�������5u�.��R^�&ߋ��Eb�U��u_%��7�r�.�8
�Y�7X�̥3�,r�N���`)/������3��iWE4\P�Wcl����h8I�J�!�jV��|;p������T����#w����=�������})�h�%��!�˴���fa������k���
���8�cZ�&���9=���\���C�J��S������I�D���$uݩb�����&�йKDK����<��z����$Q{�Qf(����wU�~�����փ�4!&&�BorI�$C!��>H��|�l�n`�]Fe蠖T����x�e�2��16Yz��Э!~�����ß2;W�-���{5�9�hjl�a�����U�A7g����nc�"@!�Ұd���C�Q�;AFz�Y��ؘ(���\����H��c.��gZ����hQ��ա�M�j|�\��t�RR�u�pV7�x�%S��5�.$�+����n����m]�|$_�	 \r�72���A��F�PE�WL~K��t	�z��T�D{Uh�}֊��<BM"��'*������З���B	#�#��օ*gj�J��;��<�<���ɑl�%g�E�\C���2g,&��B1!�C��U�c�J �Ao������i�C�N��I���B�8#�����q�أ�����!m�fjA%Ś+�z?��S�ѹ��ӒԨe:1K��]"�w+�#~)�d�q$ޤ��+=���H���eȜ3�.�@t=x�� ^�^����F���H|i�@Kҩ&g�dJf�ʡ6�/�b�4[4*��I�z���]�s��@d�[2�cv����]ޤ�l��H�O <�C
Tz�(C�4} �{�-_���Rn�P��Sa�H}�����2���f�X�<#X
��w-�]�;r�l299UB�#���U����g)W4ZW�9(��/@|K�q�i��1��Lk3�{C'����z�����=�
J�]ݼވ�t����Y�H}�9���a�C��~
΄�1ҷ����韹�c��v6Z����`()�b��C�~ �ay�q�ad���<��}�8�L4]oEoL�I��Û��o02�9 
���AMڽg��~��LK����l'���ɽv�l�O�����.e��A������{EC��������l��6�w����2�� `��=�#���L�F�Ռ��s�'�F��njh����6'{"�q{G�~��<���$�A�����eG��]W�����n�2�2��� ��t=�>��L�\�:�L�(�
�tQ�Qe���~�/Bb���Ғ�}@�3'����=�Oa�$��Q��5�{D���;��Jw�,�&hq��,ۡ�`�[Rm�W�h��Mq�ˌ�$n�Ÿ�a�ֲ�炧��bR*y�(ƛ��t%5h����=����Zs�X�q�{��;���"�O����D�>��sx���ǟ�tN��۝a{hg}!�r�2�:����H?�|�;}�s*4�H���Gw��W��:�\\u��=֎���w��(�=H-tߦ�Y0�=��fK��1�x\QTd�I>��%���Y�������)HzGF��>�%���RufS�bYJ>��*B�BI�m?�[�u�Dc�py蓻���dD�W��+��wG�`s!�������3W'"��o�vf��k#�ӊ��#l��T%�|��u�����C��u����dc�IH���o�[�K>������\�D�9խ0��G5�i�w0�M�j+^oą�ah�r
 �%ݭ�P]���]�&�뺞n�0���G��I��;͏��^��ԗA{/�^����3�F��_E�y�Y��m����{��3�߉�-o6P�(��3�[Ϥ��fX}�0^��A֔챒ԙ��5S}{t��t`� �Oww�8�d}�\d�Ai�fJ�Ϻ٪|0��� �!�]�x�̢ؐ�w���Ȭ��H����Sp��_�#*�{�R�GM6�i(�µ9�P������!����·�Ui9�Z�ׅ�S�f0h@�d?eh�#O���lV��҂H�
X��T%�+�*� ��}]��������������G	]|O$!����C��1�Ӌ����p�YHp7�3H�Q��c0��/�C�Y���J5��-l�V�5�Xbl�zy)s��DI�$r���L)ڋ'V�.��X�:��4��7��3J[��2���͓�v�rJ��s�Q곃�j Q0�ߡ��:
�"�h�#�}�0I�6p����c˼!+=?c@\r݌b4�m����x~~��1(�kzl==YVoՂ�g�g��x���B�YM���+�2��x�鑩����U�?x$%ܥ��s����+�ѩi-���a���Qs�*+��I�ˮ�cb�nH
�/G�\R>��[�$�ar	�=�|���hzd��,���t�v4�gm�&z#���`,�<	�,����{����ӌ)HyE�p�ǒ�
�z�y_�oo���,s\uƲ}�A��#1��M+ίŴ�T�����n�'����w�Gvi�F�0c�SL�r����,[^C�,�J�����j�u�- ��y`����b��'���]�%���P2���{�Rҵk�G�}c��?�<F/�}�dԮ����Ӫ (��K�)ف���5.6��"���*;����D�w�X�
س���C�j\�yh4�ԃ�G�����l\V1u�+'�Q$���3�o��1W��)7�-)�>�@Y�I%�s���x�]n��Qh�f���B�85
EQ�m���Z��u�C����k����,�f��0Z��y~��C�D�����T�2�
n4ljr�Ϣ,�h�GMs�0�Hn�P����up����� ���O�����0�UȈ�����6�>��g�9��qD�(]'c���v�7�m_ւ��$�����e	��c�Pϱ�r���
�����dF�0�ޛV�sZ����Y#��HX_A���ؾ�a��-r)ZdUm���#Y,�Ok�&*�mLj�T�[�9�A�o"O������ps�c5�41�	�R��O%^��S��y`��<�d�j��-�9"���y�Ec����T�= X,��� ������d�L�i�������;Pn�o5��t�������v��n|¸YQ�Ai^�EA1�#1�i�˕��"��p�d�I�7d�P���
q���ݐL���[Q�G�?�~�~HO<8 $j�|�B�9��(�7���<d���W����GE�aM'ڽ�}�*��� Z�Dѫ9=b��OP���+����Wg��g�JƼ�(�4�v#��s�)0-b��GX�,�9״LQ3�I�@�%�;����s�A��C=���A���1��a7�����l��
"E;ěe�Վb �&�XR�Ҫ�����J�V�|�[W��l�ANM:��z�Z����ǿ��A���@Syb-9���l|?����6��܊P�*�#�@�W>����W�.��<��Nwy�h�5��F\�)���Q��b��-�5:��,�I%����P��\� �zR��I՗C�2l@y�a��(%Gү/2*���uM#ʠ���l����$����2�����0��4:B�[-\����Bg�9^��]���$���⮼�����S��6M=f�@Eav�j퀉�8�[j��6'u�36A����w�,�l�#�ex�3��#bL}[�kW�C/E��ғ�T�R��U
7��T��8���řs�z��|�W��sjFq=F�Өn;�k�k� qC� ���2��Ԗ�����.�qd&G��@e;ٛ�Q�{���g-�EAl�@z"�uO��IM�ؙ�K��su(4N�������ATU��E�{ww�!�2b�@�U��:�aMu��q�@x�=�Q��F�J�MF?���R�����1@6�<&�R��K�ĒR�1�8k�Ʈ%c����1? �3���frC����#�P�����fg�h�J�\Lv�+ �z����p�H�P}j6��)#ڿ��v]�m�Qv��O�d"B
�
�D�r��)���k4t�`?p��=��:Bg{U�<�^M7�g�3��YB�"��^�*B��m�~�l��l��n*����G�7X$�Mӯ��|�G����K������Ϡ���mJ�[h<�P��Qatݵ��o�5N8g�Y��BJd�Z���_<��}�U$e\������:��'/Վ�J��>�~-���ߑ6ȒS�G��i�k��0��7�E�E�v8�7���(!.�˻_6$��.�$��B�L�o�h�$������ܑ���8�Sǝ����q���V,�vY}���w��|ep'�8T7���xZb	��ط�K�! b��~e�+�Q���!ER??� �{KW�0�~��}��5�@gy7����/����"�y�{>���o��=���S����t�J����j�ޞiPȿ���C ��r�%r�k�A�����`o<k�yf�
�zo��4+�5"�k��/� �	����r�u��Q�m���'��uY�a[z3J;�P"n��m���Jb0��NI�N��z����.�*�ݚ�pP�jU�2� �G?�/_�M�YDv�Ï(�c1��cC�
�N��(����� �� �T,�X�t��Y��Ӈ�\f��[�R������!,�U^��e��ZI�>酬O����<^I�V��a�����|�R��*FZ���]��}Z1��=�~�"�f�e��R�F�(�� �.'�Μˉ�H.P��m�|;�`��$�0�˕Zg�ں��%�� �2� V���T"$���~Ҧ�m�v2�(����&;W̱�tZn�R�6t�b�&L6�:���1LJ��\�Cx�cK�jX���3{M+���/��EZN�� �w�J���+�^Lj��&m�H�}�H�Bn�\V�v��_o��o�Qϴlɐօ5��5�U�Y����������m�gΒ�h6@ ���+��B�|��Njԩ�q���_=��a�m$��	d�+�R�Ke�F�T���]�{y�Vf��l����4�[>ӱ���!�̚�T��i��AF�%G1��:J3gb��O����,�Q�!��'R��n����W,��t؁H �JV����@����5��]�@�ek�F�)��!��i�DuG]���V��lT�><��'%������P;Z�<�
��!�1�X[�� ���jFTeS��spH�R�:ݳ��t<*qu�/����>j��Z`��ǧ�Ɉ����}�r8��֕ˤ�g���ʘ���w떞خ���b��9x��T�0��Iߎ�0|�b\��M'����涢���\��<�w�9}VO3��^7���5r|��E*��1�;f�׶�&���7�N4���b�~�y�B�Ѣ_t9S�t�һΗք��8�Ƨ7ݫ��h��/A�H�5n{eY��"�޷&�2��0� fw$g����#����B?T�S-98aGʁ�Zh!z�����G1L��\ا4��	((H:�F��g�t�>����ܬki2��^�.cb\ʅ� �֩D�1�9NgY�a�YAH�a�O�/��p�Xo]�]vyR�%yC��Je!"��r���y|�����fv�)����F�(�����s�/"�83�h=��3�[|a�6�,Dc4L�!���5^�֐o������>iq�%s]�n�TK	Ě�y靉uhTJ�kL�P��r���lv�9=T���÷���O� a�NI|��j��/�9T�s;�Y�j�Bi�5�N�V�GT�X/��Y<<:�)0D��T��)�m�+�!:�.�ᚰ���Y��ku��5b�IP�Ʊs����4\������=�9�Jg[_+��\LEa\����3��A�����Y�f{�,��Z�ϊ��#o����A8���FO��� No���C\wKǣM�J^_sFVͧt{�۱y�!���~�S���á��q�w��LĖ~��ӑ�;W{x���f͜m�
<h8���*�.;�x�S7�/�]f�r�nK�
�+�Q;U�,���52�fϵ3��^oG3ȉ�yY��K"�|����ꆘFF���	s%�PD�C��!^�[R�B4j>���w��G�"qn�9��@4���	_�Nq��$�6�ϰCS�d(
d�S���l	��Pl�Y-/�9:P�B��<��{e�I��Ic��a�ĉ��w��s��n�i�2^��#;][ld9�r/4nC�R]�g,���Q���H*������R�z���6lG�h&8R�s˧�����b�A~��bFZ�8bT���W��`e%ux7�a��5������rUǶuJ�z�>7�iL�e���A�bO�Ժ*S��f_���C�ʃ��4	g+�9�#o���>�PY�=BY�h���%$#Q���uc⇽R�!��RC�d��čoN.]-u���f��^0l�|��;����Љ[*7:�
7���7�=��Ŗ����?�Y_�L�*�B�N�=ͯf��t5���3���	6���F�)���c�sS->������[���Y^�g�U�1�Ӭ����.���Z��	_����f�'>a�@�*�֒�<��#�fW�Z$[B&#\�D�5��陥����"���(@�	87 �6��c�8�K�7r\�ť���c4��{uʽ3���k0�1tE���T���h�c�;M���D�[��%:AI3ƣ�#�P����GNʊ��m^;`�IYVW�wi>��6ٗ>U8��9�UpT�TFS��#=��v����bs��n���[�l
����5<�����f�b�N�����-5��@x�:XOA��H��ʹ@��r	9(��3_m��5pY��s���l������-��Cyy����[��_x�5�ƂBM7\�,/E��6�X�n�-Dc����O��<�m�1wc��rj'�:����`��7�ݿ|�"�p��kO�GK�y�տ���*��������D���W��0[�U�ߗ�����c���������y�lQ����5�)�JA���5�~�ɩeQ���I�@�,bm*��5��TBD��� ���[�͗����S-�6c�E��:e�R��6���v�ŋ��-���U�k�G�Leu
$�9�v��Y��+D�LW��	�����|��z^ ���Ј�տPa����ȃq��������m:�\�"=��uYr�8'�u�<��v`���K�3���&��+rcZjµ�,<���]&�\���d����R_��]���A�%����⨅��$�&u��/�<�j�IzQ_ч������#�%�O7�U(Rӫ3]40ə;��a�ʪ�sy��u�����ܩ������\Us;'��X+{c���c�9�4�򲂼��T���F�H��+$H��Ry��c�P�V�#�Յt����͢�a
�����\aF6�Ri��r/��ü������I����E���Ic0��i��,O^�1K �F�%/#0��������B�{t�#c.�K�8G�`t��1Y�:a�D"��U;�>8q⻮���w�H�ݛ9�*���������	�q���<8�1!����E� A]��Xj?��'6A��E� �[�#P0kL�'%?����Ma	ȃ�.-�$�j�9o�(D�E�E�C��b�<�߇�i�e{�z�)�'���m��Kǌ�����jMT�'��ҍ��9J�9£���v�������Q�=�H�q�*���(�hû�j	���F-���сBޓ=� ��Cy��5���z��6=�9���$Yz�Z5�|P���u�g��t�� G��H@B�2���^�@�?���{cq�ev��'�E�rֆ�8��J/0�|ف&�ɘ?F:R��^#�F��v�)�}0���w\�8�z{%N��c#���O��cw�rzh���ө�B�=,۹�t�^���c�������fp���X���Ҁ[L�[�Пm;��Z�\�?b�c��HS�)W֭0�p�Ea������?��8KC�J>���ܟ�Wf;�+�TU������zҔ��qƉ���F�%��C��%1�Yg����K�ɍ"{(�/�%X^�^e(ڜ6.ܥ,˄��T|7l���'h��ax	Z�TO�J( ��M���}zfF13G%��J���G��?�e��F4��EK�fW�J�w�&�(��4fW<;�n������г�I;Y���7͒��(��8rg�Ѡl�m�g9�Y%&.0�u�	 �kT����?d
kҮ������R8��ykV�	f/*�x���.��y�H�R��q=�@5	`��CQ���;�
��{hֱ�RӔxyȍA��v���l���\��CMF������w�x�2���&`��D1�V�w8y_u̅O��j���8�q�#��+;�� �:��N�}'�!����CT�՘��Ր���7~O�^��h�vo�`h��ʥO�T_,p�Jg9ފ*��%Y�Yh/s[�ɶ������C�;��,��w�I�r;9IhÒ�`dV)G�f{W5���}��!|mr�׼_�_Xo*A���%��OVUD|�t�TvX+@EAM�H�3rƀ�!���k���A�P�r�Tj��	nQm�ַ�:����M���Q��ڢ�V���x�y�����A)":a� s5;�t�Su	��P��h��5�$�4�wM0�ڴp���]H� �L�f5�dx�#kBS��Nn�o�!8�4��䲏�`��d{����ح	����mUnf�o��r�]�����2�G��+ᚫӛ��_m��ajZ�Y���x���_\�n�L�ȴ�c<-�1\ќ�'�H9m���,��n>?�eɲ	����H�Zx�I������?qX�3��iU]'�T���FM���R�C(�a�Y�)�[h���i�u���>"Ԑ���o�oc6�8���Ј'�%��x�a���"�X�ѐo�Gk2�$D�9愞���"v��?9�s0�j4l�q�*�k{����yܒTD�'��~S��f��{��;���	��Gu�o�\]�̇0~��!?����T5$<�"�뒳W;h�{7�bR�h	���|�51:�G�\G�B]�M�f��=Ǜ�D����S_�[��rd*�7��9 O�Rw��wYj��9X���@i�ln�H>���k4D�tL�&�{�/�= �zLf��P��P�~H|���2	��-�w����,]]C���+�Q�FR��yț�b�?�0u>��Ɗ��F��Ia�L��7k����xY��,m���M��j�v�ЌK�L[DZ�M�mĜ����P88��5�_9_���z~�/�n������q$m{9�B��Is�S�ۥ�8[���y�0�����L�jnܾ' D&3;<�ѯ����{rv�a������f8o{k�*�B�j���ޓe�����?q�E"�?�Ƭ���
.1�OVKn+H�� ���v�'F��ɵ�+����e�u5`�Z���D@�Q��7�υ������]�QR�︛=�a_�e�$yO�cs��Î�Z76e�~��PsHB�a��cq���9�K?�4J�PK�� f����h��V����$�Md����Ԑg:��;��(oH����Æ�����6�9�td���g�B��D����C� X��&�1�l��$�><��CX=�uau�j���'?Y���YZq?2�>��c$����5hiԘHD#�b��&I"W�G�x-��-u��򋒸	��M>�[�'�&Y��������4v���P�}���d�x�� ��Q8�����V�_7�n~���|`	�^�����k`C=�*n�����O�/��'L���7ye&����QN�ӝ:�&I��e�d��,'�H3�oס��tZ�"��Q0_�el}�0����G��qӬ�ec��#je%T.�-mVO�yҥ#N�kj�W�;����%�C29��?4�x�h�fۋx�c35�H��'��w
x�!�~����$���jMXQ�W��ps�.����|��6����A1 6���[��w�������/��wMXA��X�.�r��ͩ��A$D�M�j����!_��V�^�F6Oiq�xNA�iռ���~��!>�X$sb��F G1
��uLm�h榳!�>������?r�x�m�s�Q�s8"n՜ߝ N�1���\wm�)\��	+>p)tDS�y�Rg������5�@���D&��d:� ������$w�i�3��.�RxY�,�ҡ�����cI��^�6�vZ�.~�_�����L�<vq�5�*r]�``S�Rh,YI�ַ��7A�}Y�G�k年m��ay�b��ᥑ�{�2��͠����HF�o��>��̰z�f슺�jO1�>�$)ӯ�ğ�����ܰ���(���ѱ#�w�	�4FC�����}^5��U����倒F�l9��b�����2nOL[�o�h��Z$�ө�L�2��沮�x
�\��>��r"�^������20�_��-��. h/�����ѿ$�f��u�C�hطwayG$:�&0)���c �av�$��u�\��e�(y�.���!�����(\��#�.���|E_�6��ub�S�IϾ��y_����p�w52���Hc�4��b �J(K!�����i^@��N����h ES�� S�F+�N����]8	�P�Yz���K�X��o��/]�8�[�}y���q�IW�b]f���&�&}�كi��5�7�����=.���0�(.�%��補ʂ����0�
krWD�1�(� �M�U��W*E2�v��npYP%��J�����������:���u�h�X;��v/�mA����q5
Z"D/�W#�� 7�� gh�ߨ���տ{r���|��h����Mz^fH�{U�R7�����@b�T��HpzL��fҼ������<h�-`������U�$<d�P:�e���[O�-.�T�,K�D`��ebiGTB́Y?��U�9�r��1�/���.Ʌ���B�L�|�d	m����VXJ|��+��:�,�^�(XpZ��E>H���FB������Bʃ�o���)�>�ʭ���������se$T�Z �Q9.�w�$Es����IP�X\�Ai���>��SU7����_�TV����ZGs��a��A�U��Y7�� w�����C�Cۥ����b��Y{헤c�V�5~y����J�~�<G�!�����32�δsOwT`9�(�T�KAX5���H�S$�a���U+��x�}I
��; ��Yeē��Y�a�U���TRҘ���"�wTr�����ܟ*P����n��s�B�SP~�b�6���s��e�E �uǋevz��G�zc�'􄄷̠�k�Y�]�}�E;��G��H�����H���^���tફ�ZD@�C�2�K�������yY�R]ڪ�8Đ���#��,6#���?���LǸ����4���UP}�N�P�	�h���;���fG�.��6���@�%����s<�F�:7F�9f6>����� �++AL��M�Z�D��%�c�h�ЬRS���i���Ŝ��Q{7m?/�p��'s�����4b"����xޟ��\�|%�߻�N,�C��O+9gq`�8����'Qto�,8'@�\�& ���L� 2g�s��ڷ����I���h��dL4�L!� �=�O�[��e��<�{��s˝R2�MGЂ�����_)]�s	 ��)y��<ڙ)"(��� ٺ���=M|����	�_;s����)a��F6���qKbe	�����2gg�`��q�u�&�ib)9�/=ǀ�hڗ����+F�nqhј�~X{I�_\�[��I�n�d䳑�l�"W�f�r*V05���.�QݍѣQ���D��[Т��6�ϗ	��fd�Q�p{ڵ*��Q^�Қ�Є��#��v���}a���`�(|M�x�Q]��ܵRT���.�NTtq� @��/���?}(��7�+�]%E0�_ݎTU!����|���L���"Q�JE�������.0��7��J����������*a5��7��F�Y#r1@�s�{�S3�'�y�[�;~vX�T<��Ƨ�Vf0�D�9i+�*� *��6'�ք��*�è�,�	\�V��|H�����HF�0� �\�c�ȴE>K_(����t%�Ls�#��� ����B�
+J�/L��As�}�.�� |�`����GUۡ��tiuh{0��
X�M/!�f���B�������P�}�N)����� �H��iy�1KH�Ȍ���
X9���S�k�������L�OB�%��8k	Y9�V>9ٕ�")e׿�`�֬vti��7D��8�����������ex&�3{��KSn�:L������h���u?�acxu|c��B��dtYm�1P%z�o]p��Ѳ��#;�%'2%O�,% P�C߇NPQg���ȚD��x	�����x�hV��8�5ܘ$�K��'�c���鎁.�=�{c ���Ӗ���9�e�(b�X:��^�-�o��iW��s�����e�1{=iBsS���	 ������"�n��N	ʧ��Ƈ�w�~�����2tJ� ����Z��N�ze�e�U;�Ey^���fW���No#�qx
5i{�kiY��R���m�Muȿ���&�3�v�.��2�����fT�_ �'�: ���uښ����rV���AQƲoU{��nx�����("I� '��v&�����5�:��3aH.��/E�t� �I�\8gɧ����%~U(�")�Tٟ�j2��^~�w��6���B֘<�"��u��Leݣg8i��V���xԆ3p��C?�8y�.t���.��e�Y�� Eb��0��O���W�A�蛓ؽѨ㐭`�˕����d9���p�?G�C$�C:7{�h#�k��b�(^�H���!Z�{X��4y�	GՖd�b?<}���i���������ӥ�=Zn��hʲ��F{^��s${q����T��.��ó*R���Ԇ�(���I!�s	/�ջj����]̍�|�YE1���dK�=@���eT�,�X�kP]J�j��!R�@Q6i���=M��Y\��#��lI�?�c	�~Ӌ�г�5��L��mMq��i�Ե�E���q@�/^�#�DD�"�Гy�Y�z�8V�Ջ����vhN�����^j�x�f�>W����Z��,3K�B���L����BiVʹ�C�,9�j����)D1�������5#S����9A���r!�H��CӘ�yR�bMu�
n�D�/�8eNLD�f^S9aP+,�&�|�����Ovb�;��&��F#���_�*)��V��!��	���K-d��"n�x�ub3F�V<Um���>�Dݯ�d?��2�OhC�5�0���
@?�.1m0��"HX��lq5t��
�vnF��|��f�^Wqg�F��
���L��'$�s˚��W������;d�vf� 3 ��D7E����~�+Û�w�>B���,��H0GŻ3�*�����JMYJJrLdU��;Z���/���,�d�ʃtm���Uɍŭ�m�<�fPX��C�P(���>z�:�Cُ}��3��/�3֤sg)����!>�t��Z��m	��l�߼QԮz����g��������]����K�+�~X��24f�~��=���o���_��
�v�k��뮱���jό��*"9'���p�"�|d<�%�>Yz��؃�����pI�Vq*0dF6	W��o��r��B��b�yDw @��PƔ�DM���`����4�4�#��S:�L��W'	ʊ*���#�:ϱE��t���1<Tx�k��;��¼�I���f���^Y�oJ���y��b��^/з�N.̜>��P*�>� �F�~j(�}���Y�!��F.���kf��^�o
l�a��_�����d�4�6<)�s/�o�co�r���IҴ�*F=�4L6D��CH���^������we#ށ ��@�V���1\Awf��>o�Ep�F�Y{�7Nn�������B���&T�T;R�٢�R�4��<�N��N~�ws�U��(�;W
���0������6��M]����v�]���<���Q�uLq�_��i+�V��lV?��6�
s��9���Wl(kD���Z�\d��ɸ%{AɪTŸ�v0E�cNu����t=VV}���d�k�ڐ�Z�sc��W�����C���FI��Kǆ�AnK��Z޽׏1�UMNB�����s��dW2�*>��I�m~.��M7���r����<q 婤Σ��4 ���:|O8�ƀM�u����r�*��*4�j`e�VD=�%���Df��(��Պ���jh�Ʈ�Ø&�߱Q;K�]�4&������Q�隋�)�)}��s������뭊w�5��c�6�	�^��C�
Ѧ��3B���[�'gB�k{�-&,��Fh�1c-��c��-��o�~8���0��_JE�^����n�zw (J-���ۻ�`�tHF0�|&ԉ�)���o't0�c�Q0�IZ�J��g�-.������P#����H��`�e��,L��S?�r�QfFuz��S]"̡��P'�LMFBeMiX�J-�x��]��$���\��P�z�$��X;��W�QD1F��g0����bx���+�<`��L�=��RQA�o����7��B��ct���x�ŷ��M/�����zEN��&1�cS��ޥ�4$d #��c\XJ!�Ljΐ��e}��u�g��[e�R0�L�bnǂ2�aNxOO-�g;�S�q��3�%6b9lE�����ᓥٛW$v��Tf�uY_]�!��K�<U���F�Ә�ԑ�3'���A�'"œ6��%�m�;MC$�lPɾ?B���I<�[�5��9��<a�j{�"탵�i�i�3\W%�#��=�u=�1�e�C�>R	g��x����:d(�HՕ9H	�8�U{j������ �$��n2}:���<��f��yn	F�G�cҺ,؞�V�RF��$Hj�i/�6h�!�nr���aŉ�[*�h^%�a���e�Yz��Cu�9���QU�!z��2�U�X�-��гH��j6�6�Rxy����y T�u�@F����/��p��De�	��V�TAJ[�K�-k�Ĩֻe��Nؔ���V^�K&�	�����L\F���ߏ���p�.����Y�| d�$��,k����!IH� 8�u�H�F%�3��|�s�٨��+��lfװ�,K'G�	����������+��UY��Z/pF����5�W�"*i|[��Ϧ>�bD���L�s>>.Hf�<���C��Η+ۄ�ψ�A��bP˝&o�u��QL���^֐��q�-�|g8���`1k���Z��0z���^��$�haYt���{�$#{}�z����/�\������O�+l�
X��z��;?���*�Ͼ���ޒ�a�)��J@��Y�����џ|{��׈5x�z�f�W��7^
��1��WP��f (��=�!��=s������3MN�8�&jr��
��~6KJj��곛���ۚi�5e��Ҽ]�%!�EG������<�$������P��7�3�|1�4u�l�Y�!�9m���Tk��O���d��]�d���rRqe�O������wG�2��T�t�c@왮��"�����$���Ic�I�cɔ��oE����6L+�b�M�Ү��wb�P����9��up�>#{�y�9n��6�����f:C���ߤf��!�W=�/�W%�dZ�-&�� c}JNe��	i/w僚���!H�����b��XS�Fz5��^�c����Al�s�+�'p\'>����ͬW0կ,C�?����L��i f���Ow�-[�u���<�Vu����}��1~7,��ln��f۸��l�j��n�O��3���۪N*�<	`x(����HD���4����u/�(��H2y�&\�w�o�MP���Q�0��}aQv� G�o	��x|W��yL�� �
��2�g1n�9�ĴE����ҋ�L�r�6��_Z�����z����*6������\�O��	�iU�Ȉ_��f4���Y-��.��1��ڡtS7����������Y!�wpW�Bгp����y�h.�5�^��
Sq>���i���wxe�-�c������Z�M��~�I1M��)�R���p鮷��z�0���a|F�ef��,�x����(A�Q֛2�\��/� ���%���GY�;���P��M�͛._Q���r��q��c(�����	��IJ}�?���|<qy�I:
��R�#�#��TN�=���U�wa���Uq��'P	��!'W�����aj�.�V/�L$aF ��mt�z�� "$ރ�´�S��R^��5фY�?�k��쭹Y�@V�p��ju<��nD=�K]���Ǵmf���p�������7�I�N�ܠH(GǦ��	�Cdj��k���uu���?2�_��ϊ�B{*^�{��Ti�?r�Mv��<��u	�B��Rt��:v{]�G��h��;����d���ur��i ���C�G~�؞̧:�A��rO)����CP��� h�&���=��;��m�lX�9EV��������|z����`�Wf��|/լ ��DSvK�'[�WqB���(�MG�,�J� ����\�:*�邖[�C���x�)�u��`+P��(�7i�C�,]�C�-�ڸ��I�||8���<�<��8�J�w���l���B�,���r�p@�� ���{�@�fj�5���UX�t�a}-��4@h,��[�i�e
�}cV�9g޳�=u�%u(Y�Z�I���g=E�`���p)ĉ��NF��n�TVK��M�@I�F�;ռ7����d�ke�K�8��v��P���u���'�u��oD��h�_N<��&{*�C�Lh�&iA��A�d������0���g�;rßL�V����.�6�MAU0yx�q��Z�KZј�u_��x���ԛ�5[S�X��jf��C�
W�NS��kgcϊ�<�$��LjM��~ZE�'f���z\���*�����dJ�)'_�l\ێ����Qy�U@�g�VY=zi��A�������ˁ�%�V$�T�ƒA�����U
x�of�O5O���TS�쫎Y���Q�1D�l9nA�q��*cP���௒������K m�u7��C��6Զ�Q�e�Ce��e��Rnyן$��ı.�n�k���3t����g�a�@����q�4�]�s�O]|�Z��! �<����-L�k;��g�ȀWS%�r��G���!ύ 2w�}�>�6yx�A,	���Z�>X�����	�0��V�e��;B�Υ����E���o�(T��WK��:f�ڟF�$���O_q���3�?�3H�P�e��x���6x+����.�+�4��m�"1]�������Ǽ�D��PCK���Iui}�a�3ו���Z=I0K�t �i]z��)�¢ˑ��GX,+�8��ҜZ�]�ԛ�L�e����x����R�����d+`�U�	�K��S����;-���>��^��X[9x��"���G��l��^��ƫ��)g��-A-��:ʦ�
�Y���
y2�~h4�HM ��Q8�G"ɼ\T��%��}�!��}f:��{��!,t�Ja?1��7�J0���ɷ\z7���(�6�#ql���
�]S��\h��'�a�U��;#Z|�H��L������3��UXf���Q��k��	�vG#f�f��.OpϷC���)]+��ND���;��p� ?}���]����l�Xi�ȶEXл%#�N�@���qj��.\ʚ��n�6Ɂz�}[��bsxT}c�)Q�r�$֞�.�z�H�d.S�'�����m��Z}�\�}?X�%�S �^��+&.A�8�~u���CfP9�j*=�)�aؿ3�8�C��z�&U����N8Hz=C�W7��}Y/'Aſ��y��i�"�XKzZk�fcʲ@��� �Э�?�2`a��'�"j�c�V'�"L��6�1T��F�.��󰔑�m�RsU%"��	���F� ��hr�=�d�?d�$�opD����d������s�ej���m�"�4�N�F��1������)��e�-$��P9�����Z�v�?�%��qY��l���A�a:4������!��Wd�P~�e�x�0�-I@���w���$�G�%�",�cr.rc4�;B�d��-Y-64��~�̽m�Ҟ�t�LxY�D2����R�Q/��qsap�C_+#�C�0���7�8*�	�7���������c���l���v�iz�%�4��}��.I������X_tzL��#Ânr���{ZO�v ��h7��
-=��E�"DWw�*�T`ڂ��&�zA� {ywBm�|�h3|�������mA��n�m�$)�I�c�@�,[��
��n�/���D=��Т�e��r?L ����3�O���6���r�)�2_�L!����#�H�N	M���ur���HW�k���X�<<H���I���o�+d}�E{�~Y�����D������2�j^X�Y�сd� ��Z+�E1����P��URn�"U\no-ˊ��\��yrs
��<�g������������=�7!�q��� >���3�P����XN��C��L�ܪg�ZVy��n�z�.���:��@۔q���Ԯ�M�8lpt���~���ah�����ԣr����P\J�%y���3��G
tB���1&��k��/W��iы������aE	�l{��	���ӑ�sp���'��ꜜ�4~q\�[��S����M�8��/ ^\��ݼ���Tp�J���uq˻�E��I�#W;�D��\^R/�z�d�c�ZC���#�/�#�Y��&TݏX8}�H>����'�@(�IɿC��m m������adc���;�Mo��aHmy�XX�4�(�;I�!�C�H5���Ht�!�޵�i?w:1�S��s
��4_�肸ѳ���J�~�{>?�u��������+t2���CcPH�qN�9a(nh���Z�֘hq�JL-�o�e��F̑��;�@}ö7��[��	w<���p��=������ܹ��������1sJ�6'�˻~;�<~��]{�!��Ґ�}a=�[`�VG<���)8���?C"$
4p�Nt$���x��+{痧r=��j�!g�*̊�K�=U�ɸ[d�*0:kF�ϺS�Z�j�f��"e�%p��`����A	t%� �J\zcw҃�����"+^�ڼ
�����%�����7w��T�oިI'L���U�Z���U"A~=�J/p
R`��Pw�-�Õ�C�����Q���p�y
 �й���8����J#����X����6_ױ4{�=T�+�[*�=Y7�\��(�~��5Q��k���5��n�`/'�G?��Q B�b,~�~-+d͖~�Ezt����'>�1�p5��]�v�9"A{
s����:���@��z�������DD:��#}��a�My�s��_I��7�Y���)�]U$�+��,吕O�j��jްN�b��&�o.�A"�&m-8��v�$�ݶ�k��n(NE����g],*��ef�ͼ$3����3[��ZR/��G�1,���GD�K�aF�d�JVӎ ��-�K��A�������dkE������|/rg�[T4c�R��d�h�NGL����m�Û��B<*�]��T����pDS��\��I���0<������H��6-Ԗ �٨�����(�}?�Ȣ����f��ȡ��!?��{��>I��y���i7��b�h���-�v^�"up�<jp�5$� �� �g���P,�|f���ZR�OA��>�ǉ��8�������|������l�d0Ѩ���N�?����5V��:j|����2)�
Uro
i�ը�u��3�9�������=�F��(z+��W�`h�+��(��P��8�� �cO�/{n	�Wׁ��~L�2�&m���uH�@	�{$����o�wwu��G��0'��Cweķ�kN���1��J5����j�_��2�$b�H�z��!,ig�,�2a�!*�g��q��I3G�Yl��d_l��E���->~!����p���)�^�F��_������.�F�;d�H�::o5�8�a��X$�kW!�PD��uT�Ӝ�+���NC��� �)��f��3S�A�|Dg��:���qaǆ|5����+��g��p�	y����~���e$�H�����l#HKB�(��V�$��↜���_�j�������P����4ZS��@��ȗVF
�g��&[�-�H�{R�Lp�F!���mu��-�ڢnpӶ�
9��ʳ�u̮��1	��^#�9��	T�J+o]�5S٠
iX�[�~B�W,m�����ϓ��j|�r�j��+[p��"���M
�v��p��M�՚\�c��F`�gf�ű�(4/'�F�{&���6�)򋵦�j�5~T��+e#)���*8��.45$�?t� h�F����94��@�L��z�.C �v�*0,�J�:�k�1��-?��|>J�ZT�崬[M%/�Bcw���_�d� +�fUߛ�:���p���T����n}���~����YNAV�3&���Zu��%��=����|ĸh(���3�˃T��jA�c���&ڏnD�q��2:�=����s��r;;*6#�u���q̥��_�xO�A+9�]U�-H�^�"���gk�1pC#)���>C����'����zg{����_�(`�6%���mkN�R&}S� �)U���������*���3�|.:Y��(���Ao����)����>������D�KƆBh˖ID[�6	TC�AD��h����W]�:�q��0u�O]�bt�,��{�֬x�ս�GZ��Q�$�u%5�p�^��$~h�נzc�k��0��Y��� �{C�*X?o��G/j�#��?�_����wb�g��
��?��ɵ�����%�RW�Ut�e�+3��ޘ
����9����}�i}�ÔҀ����rX�x���6ǝ@�� �!N��r�������3ŧNl�$��Kб7��|�
�̬��������JZ���޼�\!����=��+ $��9�T�MuJ<�f
���i�ͳ^�d�@f*���x�#���0UKCS��GU���%Q�B�'��+^����H�<����ˉ1�FTb���~���*ਖnv^wy�K%���-(s_���s^�����x`."g��ʔ8l�|#�.HҌr��⇺>�}���D���H�53{���{;�4�X7Lnew�j��8kI#��,��Zssp�M�v��J%FLv�/6���rm������R��Z�u�T������Tj��p��ܫ�x�1}��m�&Z �vV{K����=�K��̍' H�&Ƴs�5r!���ݷbFF&ğ�EEYF�
�8�ɏz�ʑK'��=;��E�J���ƨ�y��R�dr�
�{5�:n���<X��r��8�D�O�ʣ�\�J��%m��q��) ]'jy�{ݜ2D��f�o��ٹ_!��a�3���Y-=>���>R���t���=]�%�xѯh���Xb���NI�4r���W�ؑh��c�dn��|�k��8��6`B~�pJ�%��Ix��߹��B^��X�%������k��V�u�?")���	C[R/�lLo�eًm�{���x
\(�>|2��OG��
�C�P��@q��O!)|���o-��M�m
n�iV5ȭ��o���8e�IǕ��oJx����.Hz[�VC����dQD�pǼvF9]�!A�~ĨgaD_)��Ǳ���w�0[����i�؁�7���Q)���S�U7mx�{�jI����ePZڏ�SbЉe�$��� <$Q=v��� ��?�P�}7A�����Z-�>��m{:�ۏ��*�d4�s���Hp�K:E\	�~��x
o!2 �^�AՓtzx�篸B�7�K����Wp�Z���m ����.�a�d�S˻�!��.��Ө�Vx5P^U��RN�Ĕ=�q����em�FIf��wבr�!fa��ݑ=�g؃2cLh�#�N~��Y[0���#��C��39�|�+����=~��G�ZgTa�$�>��y������K]�)�4؀URKI�� N|7�
�����/4�@,j�o�O�."��cG�h/p�_�u��29������u�1����cXv�W�h�&��~{�_m�����.bU"�m%I���a��:�l��g�M���9��]�������x�n�ͱ�&d��R$d/q=�1W��ؒa,rʝ���Bp{�8���.)�v�˩���M���&��s8��`�LY�s{���w�\�����ֱ�D[�E<��Cĳ[]��a�5��`ګF�Td��/3�'I��������"y�&up��X�� o{�E�݁1���O"�ȵ�~D��$ď�"=ۈ�ʜ�g������0-�z^�G9�d�Nr��5�@�FSW�گ�B!��r�zt�$jw�uT \ܳ+rÃ݋p��n�d|���O��#q�Ե����(EA�I�a��C�d϶`��f���1+�$�{ىu�Jɦ�I�:x����ǣ�̟0lpg�݄I�à�S5�wc�Y�U�&�5�+�j�+�4�N	MTg0r�&6/�	��[�>����U��X�Z$B��Gq��N@���l��	�j���_�7Z@��([��-�=r���BNV�/wn��)�^��W���[P���q%�8�k�������0�PH�]�� ˈ4��\����oj�#�;&�����πw90ly����%ky@���eÒ�hu��
-�0�	�#�=9/�d�cHp�e��~�baba+�&Vv�;���aO[���SA.��x��TH�oy9W�7r�R��j�e2<��E��N�#+-8on_����I��DƶF�(1�X.�L���2m��I�Ǜ�3�\�� �R�b�l�]�;���n�Ñf�7�4����&+\����&��}i�Š��p��*�	A���	���|R��ev7��])�oi��	gc0V�.72�\s�E���&�/H�M�Va���Z�g�SWnL��@��@����~a2��ޝS@�0�ỻU<4����%�3�H5����P��M>�@���z�ocF��9�7Ԃ͗�{2��z`W�q��TpG�RMO�n�Q�%���p�Vr�]�Y�����浞�J�a�m�:��4q����Oj˄�D.����U�������ۯ�&<�
 ��\W�w�o�>��(��ƿ�~6�i��vQ��e#����8C{Ƿ����ע��ՙ!?��Nˋ1��Mf�[�ܪ�r�2�_|�+YƋ���wC�=��^ź�~�p��/T]l��Xw��6�x��%fvBa�����aw9Ŝ�
ԏۡ�u,@>�ŋ��`JD���ܿ����Z�K���`�3	�bn��ap���Qv��w���rVQ�QE6�qA��GDFJ�4)ԗ֒��zC�K���f���3;@�珙6(������|�y��5�d3��4F{҆惧v{Q��c�C�g5;����CY��K��Γ_I��K��0� E"�s{^��uu�{�/IӮլ�]pK~��o���,5�9U�-NMo�Ĳ$��|�G��n�8'�p���Eg��U	�_
c�~v��"d��fs�I��۪��s˂�d4rUD�Ɣ��S��Ø�1ޏ��M��U�66��Ȳ�le6������($��a�D�fj��)OW�q�0`,&�����:X\��I{���/	��Ŭ�t��0�bp� ���}ZQ��Kݜ��k��� *����)���k�'V��/ Hp��=	��l'��b����
n�.$Z��e��B�ӽ�?\�@�L7��v�8N��9���m�
w��d����(��)�n+��r�~��aEa��m4���	����N8J8����������OG����3�m(~���|��sq�=�}�b@Ս�!�`�D�Ϧ�"Wp.���MRS1l��<�3�V25��������+��~h�6t˝��*r({��W�bh��l�a��uTД".��M�c�Ex����Y�M��4��X�X\�wli85=(#v���V�-z���;V�Gj�s����E�U�n���ȡwݔ�H�ɞqt{��n�֭������L�]��� A���P\��}>�,��k6�9�ݥ��v���o<)�g���>�T�(�K Պq'��� {�Y'�t~�z֓wPV�M=��PU��Χ�0ۀU�+ܽ���9}ٜ"eo������)�F���Η��ϛ���	�<]�=�k<P�������.y6�ސb�v8r�ޒ��bu������N$���#�}�������x�P�!9��!�o6@D}��縫C#�A��s��V��A�P��ÙC���߲}�<>g�+��b��P�<�s�N�+Ht���؄1�|��Ń�+m��ZX$�=N�˪S�>:	eȽ�+��|���
:���8�yS]��%���R��t�e����Զ�|x�W`�l;��s�_0c����K5whK��������@��_�#�s@,����d-2�7bs]�T��`����]�8��T�l\S�����s����]�
��|A�H�p�;|�gk&�@W�?��W��(3�������k/���Y&�)��D���Q�4!�WLZ��V!log�I�����٪����wSq)s�Uow�@��.��|/4�`�?"�|��
�&����^��垧M�Ҋ���0}���q�{()�GI���7({K��W4�Y�'�M����?U�L���փ"S�k�T�n{y&�ka���&ws ����qԱ9D� �R�"�Ez*ł���^�n�)��Y&3m&�g���T�b��(�t!�x#z�֕R#[I��i�3
�܆�2e$I�䌏^n>?ϟ�H���p�뭖1�W���~�>���ǥp�k�ǣ���$"��u����8�vn{\�$ٟ����M�\���2]�)4���V���yg�L&��g�E,���G ������C�$W֐O3�݌%����2��l�T��G_�(C���Aˡ��nq�*�?���z�Y�u��1��
����@ixB�F� "g��a8G�jO��t^(�.���߬cK��'��2&�x_��Z_��Ɵ�=��do#��v����c�]w��V�s6ڌ������/:h���w(R����Z�|�{�E�uf��3��T����b}��д����/ d���'�s]m4��,�����M�xu�C�7Sd
�d`���Gm|ʡh�P�E?>]�`큓�uNcY�=\��&Sc19Mg�}��S_���Ha�t̰R�ڤ���R��vij�7�Y�ےd�E�J_��y���w�<�%��v�pQ��P����0{���*J��*��RU�__ܱQB�S}���^�wϼo��Zz2�2��� ]�W=���eBg�[WQ�%�lv�^�Q1K��g�$�,�d#�!��lk�E��"l|��a�F#'�٨���F��=D�*2�g�l謓&����{]Km����ȭ��i�-��O�w�"->�:�!y[
<G|��������D��<J��sJ�V��9�D�ͨ���*˪׮�k�qW���ԦB{o�=3� �`I#�L��<p^�![3�̢7P���{5@�w�ѭ �@�{�m�|��\"�u.%H��i�;����l0@���6�}��9��K2��%@ݪO1���t�#;�|�.	��j�h��t�
@���M�F"���\� �4ZN��⸘��)jꏫ%�W;m�\g=&�EI��?��W������*��'2�
��#�p���m�Q>R�+��ys��'`:�~�狤â��T��s<���(���5U�fqI"S����Z�k{A~��U��	'�8󚼥���v6;>Y񒠧3��[WSɤ�8�(���c�Qj�?b@%7+���sA�bb4Ξ��߬�9_�����6*ԧX�_��{�7��u��wf��;N�{��Wy��%�c{yNԑf�}�-��R��^�&�!Ӆ~���wsnL���z�8���;�_ͧSv;�U���s^��89������ކ6i��N6��c"�#��F�������M�����'���8������lO�OV/�^�Ǘ_6���-� ����u��T�u3]4<��R쓒H��+=���,��B���W��]�M����#1�<h��VJ%!�d d��MX�� �����K��wK���BC
ލ�Ѕ:��~������0f��?~7�-��*�NX1�8Q��4��/�����!VQ/ncV��v�N�Y��q�w!�=������hX��:����?��E� _�������Yo2�t�M
�3�\JM�^D9>R=0�Y��{fc�=��%8�����G�������AKJ��ض߰�Em5��pz˽�|�����]%��a):.�r�x!��<j��چK�D��d.���>���QKUL�p�U}q��V%eҲ![�O4�xА:��M�dn$p�6*�ic#2��RV�g!D���y�N��g�O �����^�V�}<ڵ�go+�j��4�i͛�;W�tJH���|����q�I| �x�w�<��׹���^w�����2��.>�p��&5�5��Ӿpm+�kE�R���?o����I�3Il;#~X�Q���^f�h��E�q"c�Be��`9��ȗIi�H�ܳ�;U��pO��رHH�����2���F=�	�a"�|��ߧ"'�7�t,�N!�����L�t/oW�N�Vpd��cY?�~�{����b��lZ�3	�W0�^��՝��k�:KÞ^(5��,��"�e��{
  �w � �#ꂛ7���4Oq�W��O���P����㕼��ٿ�J}ࡄX���µ ��_���|���u5)j^	�z,3�s��Ie)j��0�V �dj��g`w��ܮZ�R%�)�����F����m��b �Yڐ�2������o؜�vK���es�y�Q<�B��C�D����z^��ǹ�#nM�E�8�pZ�b@�*,нo�Ll�5��lˁK��ex
��'i�PZ���?' /�ai�3C��o�q�,��G���3X5#��j�v����y�Ii�'�r��ȶ�0���bdW#^VD��9�6l��~��9������Z�R�}���̲��F�������U�%��'- KHw+[��jm:�#\��c-I���`(�7�BTٷȤ����N��:�_a���T��_N�O�x%�\2���O,gP�;n�~uQMK5z���/:���H�3��XӁ(�ż�}�nR/}	H-�
4I\r^|��q�YDk��X�@�DӇq���}o�'H�~)RLo�������ag�x[=u�8[���:�\�����8a���n����¾�Y�a��Q��b�iԦ8�G�A7H�C�'��,����ϲ^)��Vyw	I�aC�i.[R�D�:�=�x���1�c���G��UJ��#�m������|d*��u�B�R�3��5��g���f�p��m7��,�CV���f�׫i�E��A�O�֟�S7�B���lҽ!,�R#�������ǘ�D,���xo9��
�Y�m��=�\�Vt���P8��p�X'�n�9���7��3�R[�IfJ��p�ձ��X�~�.р_�	�-���g%"Ce�"߉����.����}�E��|���o 4ߕdC�bmO�5�L�_��VE�O���[r�<�V��O����_3��*h�[�]Ru����̮�6_JH��^c�'�F���˿���+E��_C���u�e����4������8�Ջ�v�N�����A��,�P�E@��W��I���Z�b$����ל���M����3ms�A!�����	]$�E��\�AUynt�2Q����^Z�()))r,"��R@�j��j�ꚉ6�oq�e|�`�O�郧C�L<c$JT�Y(B� )&c7�ÇS�Q�T�Z� ���PX��3vX�[[t�z�}]!���O��m ��Bx�~Y�m�HY�.��2�< Ռ�d�tF ]S!2��Y��~��2��1��S��'�"wD��w8!яA.�;����j�� B�pR����a��b/�ɑ�?���4h�'�>���O�o��ct�L����	����&ͤ�� ��:'�j*>q�6GѼqN����EK ��|���-
���4��<`fA��b��C���0��`n��w��v1��:z%5�J�j���'9����{Z LZ%B�q��FT ��GdZ���t'N�GLV�UY���v=V�-�NoڥD��D��� 
�?Θ��V '�MS�d2^���3�AG4����s,��y��!��_tniۆ)
�}����,}"� ��ƽר�X(�6��C��T�05�ˊ��$�>LUf�VZ�1�+8��K�&�: 9|�����^V�o�Tep[uK��,���6 ����s:�I&��}\��?Z֠,)���$x�Q���Y��*{�cu�m���PQ�dj5�{%bP1���)(ǖ���W�Nc�XD�[��cx5L��u��=̽Gý��;��	2Cy��pv6�%,N�ӘM���*6W�'�.�Ή�V�-\Z8*W����	���i��a]q�18����/`3<&�(xd�&֋�'!߆��~C���e�?��19S�*='vpұL�&���Q�;}��F�t��K�f�f�AE�P��
�[[g�V@���.e��ی,�]P)�;�ٱ4��xG3v�O��y׫��\.��1�
*�X�L�u%:Ia�ή@`�����m�����XfrU������V��^�Bp�L��֋;�����s�2�ϥ���8ozV6˂���m������Q҇h���"|3�`�,:����<�:g{�>�Ƒ�Au�H�#e���j��Y�ӆX����J��q_����Q�.H����T�\*|C?{!��qu����4.�L_}g�P(�����&�<�QZ�	�7'(\<Ԏ��6Xj7tbF~��
�Y���m��V�����3�ODN����Ɇ[�xh��'$���ڡ6/�V�5oXo�}>	�p
���{���7�3�D@.Y��f�ΐ���']ӯ����}E^$�P���Im���"x�l�Hy#����3m����A���@E?�[��̒�"aG!(Nh�PC�uG����/[bH,���!��%h8��v�;���� ��_ᑏ�h�y����1A�8k�ޯFj�F����{�O��y;wc�y%���$0DN�×Kt*쎔���!�2fU�a0��;C���6������o��>Q����<��:;�� �ٔx���8y����. y�p�aF�����c�9{�{/�(\��N����5���e��O�D�;�P�b^
L��ד�w��{�z�����O�"���d/?��,[��� ӓ�7��<�?��|���9!�x��ꢘ��\=요)>mU$�LY���r�JNo;���U7�i!.���J�s�k�0/f��G��+ �5����(��Sa]�9�l)B	��������\7��O�G��~��j]2��R��@D��UP���+����"�ӌŇ״'�mN�j���b��iK؃����g Ud
4$�Z�K �L�8wfS�X�&|��*�\�ۋ�f~�K�ؒ��),����^���n���w1�R��`$#�/�~=��b�Z�:>��\�����<$<����<�/w�r1����"��cR�!����J�{�$�$�kRi�%���yI�dd�ŉt�a�`���g�*��4��~u��#�;�-�ev%o�����j�R�������H�7k	䆰j����r	[�߉�mǒN���k�KT�D����Z�P�,�G�,ݻ�r������8#(<u&�}v]]��Z7-��|	�>[�H���GU�nY�
r����͢, �G�5��}V�X�	Q�
\}��6^����A\5Zx�{�pʅ�d:�����K�&gX�v�`�u�%YV~u��V�٢ɛ���1���t����s�@/0��g����L�v]�ۍ1�g2�$qe	o/�fU'D�Mu~9�b&�4�1-S��a���>�n�B�	.D�ܛ�%�X5f�j`p��=*���M��Co	���ɸ�����yjg���#QsD"[����ȩ��r(�*&�?c��:we4h�'VQa{�����ϥ����s���T��<�j�gv>�K�q,�lM�叴y3��5�k4�`�ߤ���eEc�+�_�cS���'{Yt���%�Q��P�2z�������yH6L8��(���(�@�,����x�+�z��:ۍ^�(����*P)%�w�72ϩ��K�0��f��Ցzh��#郅����g��WOTQ+}�Pgt��8�\�:y���n*�*��Շde�{Ω�+�
ݍ6M� �������13�'7b}�:h}å�Q����<s��+g�5��s�!���y�d9@l���}�A��-$�n�w�k�I�(
��:��+����X5���c}�a�+sA	P�z�T��*�A�,0'W|�*�#��h��C�.-�&�hQ�O�S ��q��+1��b������K���1O��ͭH�݈-�)�G2\�΍�/�)�v<IX���=���ȗ��/S���{��%���pk����4+�dW��D<�s���-���K��3���*���h�Z3N#�z�;�/8B{)��_C��N�LV��^R��V#��v�rz%��ӦH�Kc8VۡC~�0�M#1fO y�q14�A��	��r�l�j[�~q8�b����ƿ���g��@�	Fb(��Z�Hm�5ᷡ���W�R_��O���E�H���C���uk*Qڊ�.���&c�S�g��~��+�	s4��[�y�>�>b'�-<��n�I��v��)Mǲ�ݕ�4�i�W�s�ɓ�;���G��#���ɺ+2P(�c{���J8�Z���ּz�JwET�����O��4����B����9��[N�t�'MS�B!�b)��jw������{Qu��|BB�[��@��.3�m*��mi�;�s�NxO�_!��}�퉷��NiaH�����go���$�V�j�K�����7]7C��|�v{��Ò��ԕ���%N���O�.�3������x�M	֯L�<��:�M8r4�w%�<��(h�5P�HA����IbԀ�4
yE�׋"<Pi{��j;�d;��:p�JMr���bzw}���VN���<�2^p��}�ˆ^x� ��^�*�im�����p�M��-�������H��Щ�~��ٹ�0e-[g7�ֻ
�*�Y��1f-�)�)��+�:0|�J��Y�����~��D��n��WAXa��P�߸It��;���闒Ȅ�h�k���gE(�k.���V�w2Z9�4Q��ZIH����v�)��l���8ʡ�Fm��.4�$|��3r����]
������y���L�>�swj��Kj�������Ia��n���ݼ���΁���Kx��(��Qj=�>H����LIJ����q��s�|��a��M9��>y�	Y��Z�#!��L�"dXT��T���Z̵�㍅����]�L�!:�	nm\jJp.ӃW�Q��{�=u�cm���:V������T��Ȝ�*3��M���j����'&��򁴩E�*�����r?M�Ԗf����?��j�������l,���Z�;jo�Rΐ3�ԟ猟Z&�=;n�����k��	���A�:�[�Z�$�,�U/q8qBL#�L���¢��j���7���5�L {�ނn:Y�*��^B�mKE�p�>;j$�η�>Cv��x�x�)��,U���Փ��ӻl|y2M.n�k��2B����ჼ���w�;:mp��"���u����	�Ce��J�b'g���mJ�H�@P���}�=�~�N
Ȯs��nm�5m�^ ��3r04������5����7��V*�j27���{{}���0#c>���C;���yxx͈F��������hwn����v)�R���9�5��q��2UF��-�D &��XG�l8B=���ƃ�Q0���~����"(T=7h.C�uq�0<��N��J[��i���i�M#�D]��A�@ь�i�	�щ5�9&��+l���LHr�N�7l�jB�<S$x=t��q��*)�s�{u���yC����MW��I�|'?�z�r,7D�S<�G��e->�щC�`;_����D�-:@�V� 'b	{ ��[����E���^�ĳ����CR���`~ֻ�~뀾��N�5}6zujk�-�@NT�1�oTHe`�ޑ�)��3��C�+�ٝ���F!f�����`+pfn�*hE�V5�O&)�4�����7��o������1�l�Nm�M�Ɓ:N���q�1)���Fo�l~r&yqN,h�8����B��x����u�"�_�	;�҂v��f4����Rб��*����0|D�e�O��)Au�D]f�>����݀�$��L� =O����x>M�E�:�Rk�LN�K^��0���F��W��|�j�E%F=��''�s�Ǭ{��bk�1$-��VҐ_u�[�\S6��ucr�lnz�՚�~Y��.�JB������:��lUy-C�K��N/_>����Xh�$�Ȑ�
���ޘ���?)����*/�� e�٤��a�W��� }ԑ:q}��%0��)���q�{��)sCZ2ּ�$���$u�P��>�h$
���k^2�G׽�} ��P��X[�M�oiռ�Y:D��N�a>��ZY�;�N׺�G��`'����,!��8����q�?e�!���:y��3 h�yS�(�V�m�JB[=x|�l��4kE���'9i:���LW>2hcؤM�e�NP��:��sJ	��+٥A����R{�>V�� n�8 udr�>��2!@�X�PMQ��^қa;���ϩGkט�CYMH]���v<���A���Ε��y��'�R'V������Wzj���4��?���e�����S*��#;1�<���]͢�T$QǦ.��6�(=�<��H�e�_5|�F0��	��R4��)�d/��������k��$�"��f/�`$��c=e!�)�ɝ?��M�q��u�b��%�\�P�o��{41��������ɇZ"g�륷�T�*�!��X4�q�� ��
z�g	�~��5a�g�yg��������N�-���5T����	�<��φ�4z�Mn���cߍ�d<D'ڋ�1�wE��
V���!7ޅ�D��P|	�2\�,��6���]e��t��f۪�!
F>�W�Oҵ-+��~�d�IE�A��f5�	�n5�k�ń�%<��E�3VP�����~¬�#jߊ)�=�B�&�gF)/`V��u�w�[c�,f���OZ�l���b��u҇ٯ:޹�G���bm�|3�)�m=-p�1L3z��$�$��k��G�%�!H��= g����#��UU�\�"
~ϑ����Uc�h�E������;��n�����,Z����ڽ4#l�f4Gخϻș��a�g�i��3XȽ}��^��G ��c��ځ���l#���D[n׵!)� �6�\�S�N3�;�h:���r/oJ-����{�j޴ƺ�a\���D��Cz���i:��Fg����&g]����i�l�ur��q�]��F�����sy#o� :�=`*�]�2�_(��
�O�pK}��Im-����ADͨg,�	jU��_S��������߲�]�@�C? G�έ�9���ߵ�>���@�<:�A�[�EZ�In!}�t����q��^'����jßէ_\",;{�oj�dرچt@Ŏ� H�ؐɸ Ai2��7|w�]dj�HR��w&�LE��{��w�_�Z��تUH��N�W��6�t��)u� p6d-���"M�p�k�|�<{$(�CQ��/�O|���e����<�����s]��>�LE��ʊ,�d:�+zؐu�7�y�3<���'�.�/A.a����@��)R�?<���j��߾ �q{4D$��O ����յ���2�r�B,NG�D������ZQ+�������`�^�z�o���ZI�9�c+>�x�Zk"l����Ot�_�ܩd>�M�nh�l#��'i��۪6�EU(��H�t!�s�v��d�+�O��_{��R_� ���>[�f,�y�S�C��u琏��H�w��>gj4����:.d�[���P7oj�)����y7��i���}Z�F�,%���%���:��EY�Մ����X!�* MS��)J��SLn����T;El	�C��U<?�h�����@��W�3w��+���)!����^E�'ĔbP��Ju�t��,�!�k�5����t�|� ��g����D�G
A��-RP�^d�qI��7O�0iD-��zZ������_	 �Yaƹ-n5p���I�>5PF��(�փ��|��ѡ/��َ#G�5����NYh�h�O�OᲡ ���2�);�=�FJ+�a�ch�T���9A���K�o�R�eo4�ʣ�^4%���-�=z��_%�6P)���['����A���@p)z������w����Cs��7������H00��yP`�>:�!8m>"5�dz9������ɾ�x%7��|�Nnzqޤ<��e.������%�`�@� 82Jh*6�c{gU�q 8�h�6Y��n�񹟞�A}�>�v�!i}7P���l �`��l�;�!h�m(�o}
����*�f�N��XAȕ^g��]���ff�����r����&��∊ݹ���r�UX@�܎��C��g��Z<Wp8dơ����]X�&��_��Ab3uGnM�)D���t!��0ۨ�����l̓2�є΋�l'�&��f^e�et�&5�4ߪu��;�\��z��ه+������Lf�X4����|B\�N��ǌ�yT���$*���&�7Zk�0���o�����MC��IR�2��
��P�M��g"��k�̀n@�:k�3~?�[�:R>�N�m�;�a
����-�$ɴg��y�?�>w�K����t��xg�g~\[����Cgf�����S�i���=��dl*��k��	��k�@;�y^��A �Y�y	eo�Ð��7:��ޢD�nw�~* �M�,�ۤ�`������[� �Weі�p���r�o�-9�5*�!Z�^��M��GF���>���:�����㜚�0W�+s�>!vzFXM?7\����G�Ǆ�ˉ�*�������9C���T��]��<ϭ���ڑƂ��v=���W�'����X85i�����Q_x��j	\�f��In�B�1�NBxD�*��@ο�xd����_O�
t��L����Ӱ*�П(���jJE $�mG�����������{uv<�����[܄�ugM��5�{�ل���9�F�ץ�UrP7�	���~}*��@7ݒ" Jf���2��'T��̏��M�
�=�l~c�*����dVwp*G� ��,�5b�X���!ٕ��\�d?�&�{���%�22�����ޯ���5��jf�
���Q���z�5�&����3S5��ut!s�׼�O���(�F��?����;��K"�L�a'C{>^���9���nB�?��'$��0���cZ҄�"��Bo8�a�~=�1H!������Ĉ�j��>��AD
��l+�0�]$����bR++;���k7�dM��ʪ��x��"�m��\�.�W�mC-A�ʄ�w,�H�� ��Z�����l���!/��Ut�V?�{ZuIyp;*�	>�����;��Wh�Ō���~j"�;�;��-Lu�+�l+���я��k�����D���#��K�ق�&���(^�7,z^hB�H0&%z?�
�im��7ܡ��$8����KN����l��t2=b���D���;���No	�Z�6��派��MX��t�j�sYi�tɲ'�Xhq&�=�̾����><5fT�7t�( 
����Ӯ�r�(���n�h�Ǘ�Ĩ� �4z;��%l5~qp�(��2#.Y7�XP���Eu�C(kR��A��#&���ʢjP�Bx�/}:��;���@vl.��4��U��j,[�Sq⢆��m�f,�Ql�U�|�e��9�}ď�:8��G��fQ��f�/R١AiEL&�ys:���Z̃ L�M�)�	�~�/[�/ �C���+�]#L1 ��`M�� �m\��@�k�ݛ�e���]��{	�$���:1b[Y Ne��o���˹��"���hQ`��i��^`W,@d�=g���������%})&���H9��>@\��+��J̌�I�j.+.��e�V����^�fQ?ԫ�J�t*�0�ʉ����n8=���1�������}t����y|�dJ�J)��dhW��j���G�.�i�Q�y��nO����K��:�,&�O@�$�~$���):�2o]֎�H��&P�z�:��2M�F y��r~"PU�?��ꍇo�%TJ?r�*pf4q]�7��ym�����5+�np���v1V��8�Xjb�&6{���e����c��f��.�Ko�w��8n��o�jd��(�{y(Bݣ!h���S¯��8҉7\� �貳�Á"]-���m���dr��t'�&h���ۅy!�� �T6 jc���?�&6i�%q�}"��@tJ;�p������`t��J��(ʞA"��<�i����ti��H�ح�	��XQ�籭��v�3gXc����3��ŉ���K�d�@���B�f�)L5i�����]p�}���:���cK��BzDCAt虷O�H��'>���=u�x a�֓n�� r�dѢa���G������wn{��f�P�.E�Б�F�`_r�꧸[��\��m0~��
�K��~\0����݄�ApI�.@�{D���♤h�6�a�3�O
�n:��#��eh��7���#���Yf�,~�Q9>B��+%ax�믤;�C=݆b#~ьŽ��� QۘFkMZ7_X�Fy�y���+�/���PX�Ķf�I�K���#!׀�|Wv�˫��њ!��/��%��w6���+BTq�R�_j=��xk�I-)s= r���+�ĝ���:��$���~�l�������!Gͫ�*�-�e?=�jﲮo��<w�y����a{w�*��k�� ���Lj�n���N��fW��@��Ut��"Z��*��eF5+��t�y+%ቤj8;z�֖��~��~�/k~*��49�[�8cM�_�sen� s���n*>�c�2��#��BE���
�)'E8*�io����2���Pп3�"e���B�9;�c:A�E�l� 2B��I���r�A����eq�/�U��Ϥ��8V���d�Ǘv����d�"�C��N������bm!�S �����;@�M�.d�\�-3o׹�����nԚ��U-���7>G��
2�j�Dn#��_j��a�L$O8�#���Upj����u+��(��PNwZ���Im�$$x���K�&t(�ʣ\�zgA�[?:���0���2fu��DO�k_��_�����N��O��8����7����#M"=�z6ID~W�� �^n:lJ���t�M�|��v��M��w�^��"XU�u��Tُ�Z<C�3</P����NF~0:O�6�=8PF��,n��5H�h�P~��@����)�u���L�Ӂ9A��z	m2��k�3��b��].!�&/����)��֪���� �/�?paF(n��u�f��lﷄi�q�)G�듁/�P(0u��:ŕ_F햶�.w6�>Β����̊�"n�
�[��()%��ov�E��6�Չ|Xѧ�V��4U��UG#@���Yx��2��N��w�ʲ��?!�a�Qk�I����qj��nBD߀o�������`~B�m�F|!���;l7�t=qYLԒ ��&�ZR�ȱ��ms�C�%2E��-,ڟ\%�$�&����\��V7&�ѣR8��]Zw$keVƕ��k� ��]�C��,J�u�K�� ���\�)�.n4+e��M.A߷�0����A�cX4�����)0��#L�A~����߾��%{p���֖�Gx�r��k��vT[@1��Ey�t��l����k��I�C�{O&]�]�#�d���
R�e���-����!\&���Mﻋ2Lj߾�^VV0<��Nѧhɧ�̕���e	��i��zͭ�������V��ƀ�^o��(ڱ� ���-�k��OgDC�:"��W+�Kϖ�$��m���9\RA]�"mƥH�0�W��E�G�X�Zc���L���p���;�ʯ�N��{�u#i���Z�:�z�)c�!�
��j�3�Y7� 6{Z`�>�rq�m����S�([��i��?E�ͦ��v�x��.)���q����O��Ok���O%�����m��.�����V��kȫ��x\�6�0����9E��N�h�a�� �e��7�A�\T��)�}J[z��3��B+����RU��H *�"B��<������B�5Z����y�Z�Z{b,��R1�<����]tP�h={��?N�`i�N��%���-{	;;�6R�ӎ�O�$�B�XV[�l#�1uᡀ�/zr'2}Rڽ��;�r�}����Y�M����$늋N�ϽIOJ*
L�U\T}v`��|*�5`��4,U�B���*+j�u�����q��t/nm
�4��I�Ql^R��\���
5�^+s������^.|���*>P�BԔ�M&%'$��j2��4���ߊ�X��������	2~qa��H:OS��[����Bx� l;pn�q#�'+��|�l�"BՈ���I�"qT�.�e���
��X�V�]�똹�:٪bK~�t>��1��(�5��ȑ�9@A����>$�H"�����I7�	�P�����_��bw����:���k. ��6�jl5ۋ�Z}���:X�s��A��տ���>d]���z��ZWL:���̀}�V�!O-���LL��ǃ���-/���|��2g�<8��@y~��MVE��Ǒ�Ł$�#���o�m�2��!�����2~�VHکs��%?�ƃ�?�?�h�gL�Ͻ�k�$�O��qM�ŝ �-�я�U��W.�#���t�=����?���P��c=�3�M���[f������;�.qͿ3�3���w��"fH��xU�����nP��GE3ܾ��N���#+O"f��y�}�w�ތ�hA�eKR��o�l"��n�2�ܵ�R�����[LI�kv�frU'ݾ\w�g�)*4�sΓ�M��� ?�3j;i���
��5���]���ܱm��K���_O���/�,q$��0����*O.����[v�:w[�nG�4�q	�Mc�K,(��b�<��F���zзi|��
��M<�0��c˫��&~�r-E.��70yPn����( شE�7����X_�,����BLG�J��5�r4��ݱ���2�� �Cİ��0*�y!��I7@C�s��Q�)��7?����<mI�s�c�����8$@��)p6F+��Yl�K�Y~N7݊�,Sq���b���&�P�SR�0�F$N�l3�:Md���x�}hY��n;�nh�7P�#wM hd�8�Ӈ<I2�g�,ob9����ڂ���iC���]࿃ �<���l�+
���8(�Q��r��.e(�*�\B)�*bW���^��o��pm������( !��
�+Wg�v��=���"����:�R�o��A&iU�)�y�Eѳ ?-���ML8Sη5ut;��� ���?g��U�a��P�T<�'��ʺ� �z$j<<�v0<V�\��E����9BM����{D�� a��R�~)�sz|�ҼL^o�V�՟�>'Ȑ�������:�n�q�~�@H��fY��i�hB��Yn4l�-A�I�I�B�Ed{��:.6Q���<o�qd<[!���Y4*FoZ��(p?,��,��%����6�G�<�~���g���%9�r����K���,>�3=�����j�۬�	���-=x��FV_���אr�U"Ӑ�q��L�h~����_���4%᳹�=�E�͓{ek������<�7RTU�S��RD5�����@7ӲE$P��K��O�	l�`MP�؈4�	1�r�&�#.�V����srN�lD���fA�e��=Ge�����I����;��N�H�ke`J]�`o�i�XA���'�JNa��P����❪D�Y�'_C���?ƽ�Gt�(���k0�Oi�ǯ�bz�Z� U��JKDo�b����(���j��F�-�0X�3}���(���F/�/���K���D�:�˜����]���8��{6��82*[���Vk�W����b�@W5��8����6�l��::����N�nDh���e�<E��m��%��z	?7�C�ؐ#��~=U�����^���XR�������?�p�c�nIw�F�<4����d�so].�(c�>�F�ڸ���`��O��� ZV���[� �(G�@�b,
	�m���8��Gшke:U��x�(�1V�
���<g����t���Q����m�n��T6-5���.�hm�]i^o��+��0������-H8Q��أ,'�z�Nr|��K�A��43 �B�hU_A(	�dl�al*|�C���cNMdGM����}��L�W��%p?�w{��c^���J؆O�dX�h����
i,@�����
j���b�?�E�� ۉ�EH��8��hS1�*���M��(=(O��	�J*���|9����X���	�n��������.���@��=M߉�ŷ$ʩ
�����0[�ܫ���� G�-�b.#=�,aFo֒���c,������� ;�@<����G���^��v��0��N�??��{�U��fr���1_��:%$�'���A����y"�!8饌d ��胵Q�# ��'�'�O�}Ӣ��C��a�|Ƒ���8���I2a��!���|.9�����B��?�P)�!d���_��9+�5�V�=�h�s��X�{��a/	U�jQ-���B=*�A��>�p�\/8�������g,��eu|ݗ6J�����&n��煛�#gzN{r��=
Vb��;����A�D%�y��Ϸ[#��
4�{Ħ��ܝ�oR���Ƶ���e�?���B�����~��#Ѥ=X��x��_��Aś3[u� �@I��������SZ�Bc	��[�Bv�]h���O��+)��f������.^9���5��:o�ɱ�NE$B8G�~��
�����9�ХTAX��xB�<>r�C����*Qb��B^'D2�ʢ��@�ՙxšho2�٠*�C��X��+����X
�\��t�}��(ǵ�@<��nB�L.�M�.��/(税�������I���'a���^�Fđ��%qx����#��lP2ھ�7?��	��gt���d,�������&V�!y��ήː�侦�*gb+P�:�T�UY
��Tnhu+6/(�DJ��������oS6�{��K�	A�p�����6���7X���.�R���Ef���V�oI,�b��V��G=A�q-_L�4�H߳a�p��/-ck?�=c@?v��N�Gn~@?b$uh%��nQ� �׼R�T:�2��@�<��;*oV����V��;F���]S{	� ]2��E�L{u} ��x�ÖV�w���e:r4t��3������jY���2�7�g�NY���Zp���I�m�TW�H� vR8��<ֲ�����B*�h	�F�i���K�O1�\�p]�]�ew���W�����8ƃ���Ɛ_���j4�gb��J�%ǔ�l��0�@�D^:��������O�Dݏ?���-��D�3H"���R���m6��A9h�ɱ8�VH&?��V����oS�Q)�p��t�["�X'�e��x�!�R[��q̶���sQ�di4N�^��ϗ�qM78�	E� N�Ūj��Y��C�p�10�p"r�+X{��t~��V�6Y�t�Is�t�h8��3�lB3 ��kӸ��B�R�z�An�����v �)��1`;/0"��eh9��P|�^-,J��v��Pev딷>N���/#�V{�sŷz�OO���f� `Ǔ���"uY2��z�u��z�U"�&sRN1��v_2�?�^uӳH��gUِZӧ�ϻ�@��%_}ڣ�	� 8��Rr�~����y� (s�|�Ρ��w�f�8�H����v���C��bML� #�����AT��}��ǘ�����U{�)��9�-ю#���R�=kNx�lc[8�����k��,�a�vB�\n��-J'���Sw�_���E#x�[wl�ewB�"ȁ�%[`r�D�/M�^h����k��8|i���_��>���QP�{S���>�0͏�]���(r>^�����}���x�gԃ� .���O�,��7̓�.V}�!%��C�fG���W�k?|ł} <,*c�*d�*��b61NUj��E���$z�9p�T!<����r��m_j�=m�I}�I�U#<?N��se ���~��&��ô�Bt�$��:ҏ2I��"�}HI�,�b�.�R�=�Ȩ�U�UKc��������L���P@��N���Cp����>�`��0K�6��G�?]q���k�H�>�%�K=��]�D�XS�(�_-�H��U�j��>�f2�L�Oc�C���)ރ��7A>Y��,ھ�=N�x%��\�S]ɕ���:$:P�͜3`�c/�d.y�.`D;P�6�
�g$47+�3��h�zPf�6��b/2h��+�*�nZ��\�4	:��b F7�j�#o�U���/2ɲ�n�[��0I�}� "pNv��q ��4��n�?�apt�()�v��6���=���y�S4ߎ�=�����5��
�`*V5��'�SK�ruUF<���ʃ(z������F������ki��	��q�R�[�x��2�o�uH����W����k��*K��>���������z���X-D����Qޛ��D|.���f���e��ɇ��D�l)s� �ȭ�A@tn�e�D3��ty��E�����<�3A�WW�$�+,1 ��+�֙�l?�K�t�p�����$#�Bu	�K���O-�o�Rm9d�w9<L�!��7���m��]�[V��vS�,I�Z�� hj�bpK�7$�~{�:����p�:1�|��h�0��"��s,z�^���o�)4��LT|$���1?P�̣?U�?G�k���N0�%{NT�fw훶w��:�f5~�Mt��1�fB��!�����[���I}�a J�����+�[3]��Z~��yθ��.[9��b�y�y��- ��.���[��Z9d���.bb�B�u�S��ѝ)�N�(��$��K�Ж�Wk���d!����+ �v��/U�-Kȫ#4�^�k�t,����G{�zg��ߠ`�v��OaP��;_���#n�����a���t^��~c���J�eK�5UU.��8��e�`�����y{��b�y�ڄ�h�'�[~�(-kb�����������ğX��B��������.b���vq��W��j��W_M\�#z����z��(K� pq�	���SJX�J��K�PS���DU{@���aD5�^$ ���]x���6��dG��Fj�
�M���*�L�V���3r�L���Q��,����ºM�R�ڞ���c �Rxw�]e�|�OA�髏R����w[!:���\@)��ͫ�Z���C��oڞR`�k@�ڇ^���r2�y��P�ۙ�b�<���@�M*��c��(�nuf�r����s�+�V���{8[�Q��m���UpՊ˓f�;j��7������3�t@��Jĵ�!��G��ҏI� �����h�t�P��j���Z�1&�6F���b���Ü�y[�Q/Hm�F�Z
�Jau�����m�EsOBT�*֓���Q� �Q��͘Չ�~iB�ѵuz̎0��r?�/��,���}���zUJP�@[c!��g�B�yt�&�jC"WZ��#4��{w-���U=���D�/�����ͨ'Ǿ�#G���+��Z>5�K�t�N���>dx��B׆����9V�9�%�::@R	� ���V�>��;�6`���5�����ab��bvzH)p&}o�%���11�Ņ����	؏����@>p.MP_*�����0'����G������>���jv�W��x#nФ&{_� z6�ʎ'�|v�[��&"pJ�Qw�ay���b�qޗXV��`��O��}/9�C�,i[I�U�)Y��ߖ�ϟ7�������/���&3wG�L�5�Mܰ, ���������l�k�OG�i�M嫗W���=�g��Q�f�*�+��G �f�±�W,�j���P�,��W^���+�=E�+�y��ʙ���m��@�/�&dB��6�8�Q<�S���pb|cV����T����l~}|���G,�3���]� ���͵<�ru�q,�y�s6��a����
+�&��%��%�S�BXd�]�'�l�e��f��}d3ؐ�)%�1���y�'s9#QI��������k�|_�N�B�S~avy,��z�I%GD�qt�o�,����G��z"��fo��N�Wp��{&p*�?=���)l��>s����M��8������,%�bH#���Sa{θA���~�����-����8쨿H\:�N����ɦ=��!�@��(v:������u�pV
~����Z�X8��v#� i)�#���R�.����"A��d#��vlx��'�҇|��I"}	���U�������b����3����[�OG&��U�bc��
�Ո*��a_��������qG4%,<�f��dN�ڝ������x�gI|��{zA�LzL7v��,�;rV!G8�Eu�|��ҟC��/�����њM��!P3Y�n�������mxS��T�����l�G�ʦǏ��q�"���Cs���Z{L`�h�P*�L�ڔ$��H��/.{�V}i=�힐��9�@S0�-88� ��M�(p�����WK����_������1Բ3C@D�GJvS�tFL�4�hBT�6@tn#*H�.��Y}+[��/oĒeN��C�I�r1�y �(�xWj�S�I�z��-o]���<�t��8�-��#	J/�����J��tCg�0�f�i�GI��㬜���[t���a��z�$���5��JSQn!�B���yyx�y����O����-�����{��C�P���}�rC�1.��Þ������QU=��_�HY���D�M1�O��9T��+����������iI�sn&�~D�X������������l���M�<*P��}_8@�� <��&<8\��/��/���K
�k�1=1�e%�aD?f��o"5*Z[�h��@��KC�	�_߂A�O�"��E���eE4iM>��y;.t�%%ʝ��9��=�Q��M�1����ƛ患�c�bvnR�@߬�'W��Hw�I��/y����>�a�� �Vd+1ii�<�xh[�a�iɈ2��>fw���tP�8yMyؽ���U���0�����f��|S�꠬w��7�y������I�l��K.�ӆ�5�31��M_��AB�4����nƸ&�<�_�.@����DS�.���F�VA�bv,�вG�����GM����	f!�M��N�@|Z*
��"�>,Y�W�J�2S <&� #��DZ�����y���� p��K�샰7R��I˷��j�=�/:}di X��Q���Io���V�`എB�h�_� ��V -% ;D<�`t��٤���_K��*�>y�I��JF,72�ǌPɕ���y��s֪���[Ѕ�
%��X�uw�"NU��+�r�n깦�=[���Ifc�'�ߎJ+�Z��y�B]�@b������GP7��s�ܥ��Q95�YB�㑥������A��fY�<U�,�̔�p�JŦܛ�J�R,�'�k�]�⯫(�F�h�l�(���A��K]8�!m9R��*x�܃R�L�+���Wza����W�u5�$ɘ�`� *)8oX#�n��0���)�t����ի�Ǘ�ar�G��f���O�j�B�Ĝ�[������|�VFF@1�����K�3�?����Z���$		oӆu�4��zL{t�զ���95F�
dL���>�P� ������&�( վį��U�V��w:<Uq���]�T���Q�n�]��;�f����ޙ9!��f�����ؗp��;B�#da�Of�������E�%�v�}���5��ǔ�_ݙڦ��p�I�䜓�uy;
ߣ�q�[��"��;v3�Dz�:�	��^g�&@�9���C�|�}7 m*�a �e8�̢�\Ty�"`KJ��9��0�F.����oG#����_y�`��#w��� ]��PQΣ�� Tё�NViI�`�0ds��b=�(�Q��'�n:���jy�j���0~؛�'*��u�����V��K�qo��|9:�.�RN�i��D['�j�ݹC�$��е��'Bg�NoG�5{ߣ<�J��rt��'p��Qs����FMy?F��������ܺ1�l���]�{��9����__���V�Y�������2r�Sq�P(X1H�,�$�`�f��/�T��Gh�����2_�����q�@ڶs��a�ot�m�ҙ��6 gBSx\z���UA�ע��6�K�?�$q(|�1eօ�\�a�i6V�(F?Q�u=B�Pnڍa���ef��r	׃Ģn����,ٳ�fd5�#�Ȍefi.+�/���K����m���X�M���su� J��3=)�5>З	s�A�B�Δ��P$�6塸��.Q���_FϻI��3~Q�Ǘ��Y=6�eX��ܞk�Q���J�T��d�����gr]m�6��<���ip�>`���Zc7{"uoJ�u�^�U�Us(�#kB��Erehʦ�Me����SCϜ���j�A{7p�����}�y�T|��4d-�q�fڼ� ��en݅����\�Yl���¢c�T��%���r<U;�����i5p���??����'�p��܅J�0l�m4v��-C+�k�hHnnkz��%opZ�����������8��G��Pd���|�t#�ͅ��6���D����vU0~0�p�K\%|PAQ�WfuUX+2ߚ_���ʺ .��י�Ş-M-H0�����[f��#�+��{�eNg��$?�WNEDӜS+�^|X�m�?�/3�L~`:�Y�x���&n�-&�v�[���fb�6�x���ˁ�?��d��m\�n��t]�eQ*�����v,�#?�6j[@��&�{{
k�{2�<.b�0�=OUHO��tN6�?̅��z�X�h���	eK]qAaj��I!�}5�Uj� I��lv֥�R�d9 �_�a������%dy<�0|"�4E���<Qs&Wa�����@8��pס������b��zr��o���8օ�.g��̸D:n�r�,�v�gq��2"�a<�!ѼT���H�������8��{��*��)6�N�!�Ę��=r�f�Zq��N���7&[$m�\��3E���r�;����X�-�S�������gBώ�����YpM���k�0��bƀZ�b)�a8�z���c�[���Pa�a9���7�"�=�%L�_	�F�CvSTCIJ�-�v�i��І�����C�ە��7������^��tU���C�\�nEѠ��G��(מ�'���N�ԋ�e�9�<c+W09��m�لr��ӆmA��tȕ���� �/I���W"��K�g�R�e�iOe��/�Tx�����=s�Vl���(xa�qx�w���s �%_F�Szm@��ܐ�Jm2QF���7/�,�D��~�>j�]�s��"�Y����y������s$�8�}ݲ�]@��I��UωY��z
�]+�[	3}�{n�F6�L`'|�p��}��8��!,�s��
��y��LA)RL�G�Ş�XF���_?��S��Ƶ /W��[q��h2�s�@HfbU�)���VC�A�������Γ��V��kZ�TNy���:|	�
��=��; \��U�^+X6e�������%�����s`��~zL��1_+��m��s�:��r��	�"��8����YL��� uN�Q�Ӫ������L)�2|i�4u���B�%����iĎ�P�T�J���z{	���7"�s��c��_&l(8Sfb��A$o`&76�{�|e��O2��"[������������̗F=���5tR�^�Q����鍴�B�).M�����fz.����y�ܗ��)U2�>�H]�&k$�`W1ry�~�~h�������^���Z�Vܫ$�^J'��L}��^�����H&��X��1x�ߋl�G�O�����￵m��,� d��>Z��ٔN�f�LPSOgB} 7�._��1��W2�ꮿ 3P*��z�ص�2���2/ȏĖJ���x��ӖK�v{�Y�'A��c��7��`��%� �?���m=���-Y8]C�� i(
<ئ�o�X�;���rT��}<n��\l݂#�S0��;&�l�Rok�$����2����%2]��D������ #�
a#�c%4�<�����J.�=��P��oJQ�~3�����At}"D�K���fo	�Tz�Sq��!v�F�z��D�ڝh�;����9
��-�%���y�1gc��0K9���G������J��>����T����s�j�
�MV5����J��ف�7���0�-��1�
�#��M���mWiW�N�3��5��-؅�zVq��(I����l��Q/¯x�b�|�G���Ӥ7S՜tG�ێ	����ANF���"+BI�=��P!�ad��#������� X_Yslf��G��ӏ���/`¬Ai
n� Ww�?��i�
P�rɲ�,��h@h� }�[sbo�d�@ʗ�h�B���@�cC(#����$��.��<(��-��_�ᘫ�f�X��l�ǣUG��S�q��>��!��>��<Dך j�&���6�P ��t<ꈌ{L�4�%@�֣l�̃�}XJiKcJ�<�5���zF���;u�*�UhP�U�X�_�p9��!P�؝V�5:���!.��/b+z
觍�����"i�n�����8�Q]I��	zF��B�Kg�kׂ�$�a�̐��~�h���s�g�XC�s��C��u�?�e�6�Z��jx��1�:3�ގֻ�������٣�~�����2֘te��X�()>	�*䓿Hj�����>b�
h��^�5W�Əp
�4�/^���Hs5�[;�ȵ�%l]��#�$@^��v��L���Z�ۓ	F�������*���$G�XxI5g��U���e�h��-�%��b���`Cw�x��I��j�b����\'ie�"ıg�dh���k!��2��Ίe�j��浵���+@Q^�yJae���:b�BE4�f~蔋����@{��O�\ �����p���d��㲟8���	�}�[���'Z,~�6�e�0Sa?{�(��D`���D�5�c�	�3��ay���6�3��TMIqc���{�Ңp����Ҵ��J+�ˇ�`~�1�.�S�â�1��%��+�C���f��F;������Bg���*�.��e�VUw�nJ�L�{V� F�{xG�EuB��Jxy(�+���H �N쏵��Qb׮F�!����?������3�#^E�e�Jm0pH��dǓ(鶸�r��
��/���� �BM~pɛ}���#O�j���T�=�m+�'"峢�q�0Lf�oT������2���~�oh�O63F����%^��0��Vy懣�9CY�]��r��{L��e�o�a�OՈ!~��G��8��JN�z�Ly���U�n���ڤ%ן3��)�,��G�;j���.�� \N�53&W��u]�;��^��h�2SX8fL&��9�7L������U�ҍ(
�u	�ez�n�EۨQ(�i< 5�<-��:�	7@G���zO�τ0�f�QW�m��k6����g�h��������cڔ��z��k`���9Do�����QT�kF��G���4�cwfD���<�q��8�م�8�)B����ߌ�
������z_���r�\�#׭���dj4�k%�x��k�B����hOL�zVR4�lf�f��H�T^�{f��?ذ�R@-G_RL�,�"Zs�n2�rl��m,��s����.�Gs�q�^a������>�Q��*q��9O�@�9�8x�p<�x���5��:K��>��w`��R�l�[[9a��b��梁@���(�k�b�f�Q|W�N���a��B��>�i�qI����j��!(�۷~aΎ.�ʋ?�d<k����C�v��9j��U�)OrY�̔C�17(��i�ߠ�U&Ĩ��b����+;����F7�}'y��~8hWk��Y�U��m���00�Fu%����iY�e��t-8;����׀��w=���aC ����]��C�����S6R[�Ǔ�%	me���q�\T�ez#F�X&|425�g}%U�֊dܼ��T�G�K3���}��&Y��L��>����)kJ�x��3vJ��O��r.g�0�	�~k�����q5gI�Uζ�4W쉍�Wk71�L��A��+�F$I�_��9����q��8i�u����U,W���^	נ�҇���+�j�2�M�[Q%V���V3��(��x��������g����`/F�9����������%NJ�,c�0�T�'�`����v5X���W�!B�M��S@�b�t�D�ͣu�b��TLF����f�zF;�~��EsH�<�z�Ah�;������f�o��I|�:���:����$�B��G\3��̀���[�I+���2��y!v����*8<n�@��i�FT�A�9L�D��\�PB�2"�oL��%��={���,g�+ t����*'	
"��_�ͷ�_k7��9
�5\e�鯾%�zn?O$�a�[� ��`5�Q2��U?�˛���Ѐ���s�rf���<����X6��z)G/QpN�d��/1N�:�J �Mg�(�W�x�mv�'�u�H��M/�r�'/8�L&&�
��.4�?IT=��c�΁��,Q_�͗��j�(�y0�vOT��P<þu[����`Fڄ!i	��Ċp&f.d�"����Bq����3��˅�(��lo���+���,�3�/�GY���.j����3�&kO�Ż~�&!�x<Q3W*b�x?"0	4}�`qR�f6Y�/J�
;&S�h\q셨���nO}��a35� �M��[��v7�<�r�|�Y�@i	`BY�����-�'��6o2;��/s�g���ADq��aO�ߪD���occ��fO�;`�Iy�� �&+�}g%��:��P,��"���_+��v��&Y@u�oL:ck��[��F��b4-�R��龯�|�T�ۀEę��><y�0���k�s^C48�^��i3/�]�8�$L2��Mg� �74(2�H-[��.�`��-�Zk�PԚ'�=m!��΁H��e��cw�Y��:�R�8pY�g.�P
�K�y�(W��:#������<��0�T>��D	�:F�s�x1�=,�҄��!��K�6�!�>97+�l#,ۢ-	�K��樉Uo lA����;�U{E��hl��
��J��T��{-���*��-���<3�rji��3$�u������8�o���~%����շp%�Zy	��;~+9�|�����re~^�(b��ӡ�X|����VQ$���Q�\B -�oλ��o�~�=��^�h�=�n]S�2�r��O���eE@�"�WPN����%mcşuׇQ6&�h���,�H���(K��!>�~m��LGGb^Q!-�/�hkC���;k<W�g��Ȩ�������v[�˔vR�c��#�Ġ�m�3yx#�� a{-���ui@�����i�6�?�VF��P�M��`c�3>���6������c�����h��5Q���q���/���Q�����K$Z�ٔ괌T,-�{���M&�q�ce�[�-3ө����п�&a��C!$�]Q��(�f�ˋ6􈵒Vg�8��[�ʴ�E'��j8z�N��y-\*��j]��v��n�0 {=�~�x�- #^�΅i�Z���!(N���|�,.�vJ�L�T�,�4E��a�2��_?�����ZBf���^G��0M�)��c�o��p��}L��ދ%�u�9��e��i������N֛+9C/�@Ϧ����Vp\1�կ2F�W/^�|��#�h�)��b��]�s�\g �o�s�|~`q�A[��<� ��;h��x`z�f;m����I��XYo�8u��C�(z��Eb�H����w�}Xp�y��4c�V�?4��)��ʋ�T�>��xxs�Q�R�3�G���#��R����J���m�$�z���x`�X	���P�"XO�=�Yn��a��ļ���!��k��#���>Q'�7� �)���'i���O�iC5j�gؠ<�u��bC�5��Z��	�,G�C+���,�ܶ}�j���&	����d�yr��:km:u1���Ɣ��>+��\�Q��0+�k�&����ԯ�9זea���+�v��l�*Z���}��<���IzL�U�0'R a��w5��G���:aD/�G#'���u���SshI�ɇ��;�Ⲳt� ���yU�U�y('����ͻ���5-�:^�Q�����Þ�QR������1�[��Ɵ쫯j�8�+�����M�X��;>᎝�������6PKv$��E/^&� �$�lQFI�$���������zk�~�a�bmw}Q�*#�D|\�V��u�+��#_ú+d����/	 N��+�re'��ih�O��	�i�&�Yd[�-
��P��!�I�8�T%��h�a,���}x�����3V��u�8� �֢#����]>G7,��/�bYP�Cj�Z��Z�q����P���i?�_4@;R�u�1*Ĝ����}��]6�+�i:b+w��p�AꄦA�*O���%J�
����
L��BJ����%L�Rzz���3��Uj�01�%+�Z(�c�MA�%	��R(��ͫ!6�x:��B$�HO$�V����!m��y�H������Ц��_���W!��!uW��HM�C��?<�C =���ȑqI�jR�'j�mVw��5ves�];PXx�Y��u���;��H� ߎQA�XO�zOta���}�
�����"�ZT�h���ڵ�e�P�׿�^
_����d
5���x�l��`m�l�_͏���4nߟ��5�`��=bи8���)�z�,y9���j��^�P�ث��e�� ��!�ڷ(k�e��_�}�mF`��pN�K���"��A�s9�4g9꞉�w@�?��ز��e��A�Cbg�L�����T�(0�Qr���J2R7�|��ѹb������<�˘�u|�Tv�qn�)� ��x��c�+�`��������"�����*��R9���v�o�nDj��4£���:N	��?�4a �ѓ���wM#�F���w���(׃�l�4r�C!�8v�!5�s�zsʂ�Xo�A�x �U�4�ok&�YI۵�����EMJ�&�
F �����{�i�NI�H>�2�����{Q=Zjp�+��%y]/ۢ���2�9w@���5
�X��&�&@1㾂����烉T�R��<��lʩ�}�R�3��b[0��F"�H%����H�&�!�k� ��y`�u��#��t<m1��ᦁ��1��b%Kr9�{��=��͊�u���2q睂��:0�I���>�;.4���{%8#���o�:U^>�XM�ߞ����!5o������Þ�t�R���"�� � ���d`$<���w�����4�݁�G�q�����7�.Go�MC���c%���>F��?2R���+\��W1�i�����}/�\z����M�h��RO�#e˖�Xj�6���wr6��K��e����)����z.Մ^�	��.y��r�����M1����?We)k�f�[�d�hrx�D����q��N��:&���4�$��.���A��Yh�*u*h���D3���E�����K��a�wb?t$<q�.3#y�n��벯�ko�x'D\#JQ��n�҄M�0&�����+�eV2�[���2w��-R�a��:�۰_m7��)=����>i�6�@V���ooR3��1�E0FS�G3��q���0��\�R��.���B[�HBI��u���"�pq�)cNqb���>�T��;K�~N�a��!�ⷺʼ�����yn�ѣ�}�G̺xա���͉����H�50lO4+��\ӻ<�э�����W`g]Y�B{d��TO����$/��{䔷�1l2�5EԶȧ����[,�u k.?�,p ����$Y�I\F����#WG� ��ܿ0~�DW��D/O��1�`M��h���E)C�f��p�rEP2����7z�Y�v:�Ms]րY�|&�+���{Y(LLL�x�L�R��	`DV�����[O+�6�/ 1�͡o�pl��M��*�#��a�r���$,43��'���.����k�����6H��x
�擀�S-��͒�a����� "��}��?d�q[�V�2Giɸ�棤N��Kv�8S�?um�ۋ#�k��V�^'lVoV�@�C��[Y���w9��saVw[.iH��B�ZOGk�68r(D����|��<�����P-U��0�8�,�%t0o��u�o"3�0ߔ�b �`�a8��X���qJ���	!!��W��a�eM�Avt�60[X�O���ÿ���	��ٹ����������
��.�1�9f�@�-�9�beIb@�H�bW�u�eE"�.<�����s�a+G8�� ��B�*}��̖����3a����2����k�d�8��	��7/m�|f�w�J9?/6&z���a@Ͳ�go�p�j�c%������d�Li;#H+y�]%d\M��Z�Y�ҋ����e�so�x�&Y�[���]��^�(
Tyfx��NG��!2���Z��̊�BJk4I�~��4�9_$��`͕�m����͒���$�{� &��B�3��b�_�_5]"�YC�,�D|����Y��/�; �0@�C�uJ�[8i��:�I{"tɮ+.�3N��r��K-�����7���%�m�.˂|��H�KS�g�O�+�� L
�Ć�!�eo|�4�j����#,!�9�=UL��r�=�01�����KO����{��=��%��f�&�R�N����Q0Y�}�@B���c:�©<�=���ճ�i'J�!��� �G�z�:��J�dpN�n��)���͞rW���fP������v���q��Z�DX�9����9����j����O��]�/�����<����	|@i!)ID��cy���)�ĽCP>	�lsw���>��o��P�S/�Y�������hTج��Ѡ�0eOy���p�� ����3��B������f-p���0T�ms���\p��Xٖi�?Li��ݾz>��Z�S�A��Jt/@8#�6�7Ǖ J�-x%U�-A�փ����,%��:Z�
qɬk�����W�V���>��iym���,�[1YQ��x>�.�J����%��AQ�I�I�݇���p�Y�u�0���+BN��.��p\cK��w�+�N��@���b�ʃX==�R�À^�bA�H#Mc4���kkġ��j����3�fO��S]�I�c���@�{)W�*Q�˳Ăx�����N|Է��ȋ��-!\��̄��ˍ:�|���8|�#�i�o!;�?��,��{�C����h�[Rzo>b�^���Q�۫�$���y�悰�[�~�r���-���4�j��I��,���D<U��W@+�l��[��Y5�2?�3�:0�%��|o5�M�t7�}����/w*�"*�/eӶ��`��j�'�OxN�LB��Z3V��Ts_��*6Fz�$fw'F�V3�M�th[��lidRI~�豿1�<�;k���v3�5F`����O2��=ݟ����� �]F�O��|�� � �e�}�����p�w�ά�ޚ����b0]'�X8܁�8���nׅ�#�}�a�(��vp2��a%����h�	2<?��!o�v\�{;8Ӫ���]黯�Me�	�C�,���:�Ϫ�j3l.���xw3�h�%	����p:�	UD�6!���Q�#��W��� ��jE&�1�:H��LѦ
V˙���b��u�|�1^�cd���yo.[����"$#,�v�;���N��\����[�e���I�럅9��T��˭4Y�i:3�:'�@d{�,*W�r)�I��p��}�=�õ��?���3_�
'�E���0��	I7m�P��xf 32(j��M�

}��M)����C�2�TC��k��Y�A?e�G�r�ʴXv���C`���y��D\c�2!��ۅ��2��e��ҦJluzuGq�ͽN������ �2��_R~N ����!����l�&/�-�9�abf(�#��U�b9�'�<s_;.aӅ����#��@^Rw�Si�{p��${�����׷N�	ٙZ/��z��J�u�����C�*�N琑`:L�*	�{�Е�S�H�����j���#M���F�_f��|�Litz��U���*�Ӄ�]V��9]��A��IU��-*�
=Ļ���l��S������8����0�!}ˢ7{?�\,t7]X���͞X�������w�'*�6�zm~��G�d$�u��� ��4�������=��v�D���^��v_��[M�� ��Q5���M=o|S�#d\�$^�#摤;��}�����%��ehM�����i>E ���Ts8���{n�� wr�Q$�l�eY�f�31��f;���cj�m���3�	����h�9�8�o�A��4_M�\�Kni�� &CD^��a�[�̮�)�,���B)S��GY�i���5T���������M\�`��V���$�	_1i�8P�	�&��4��u��o�T�!~�����l�8E��P����d����.l�>h	�;_������R?ì7ڻމ�*b��`��bWm�H<��Z��W3P�-r�Z�U�������ux+X�"D�]��m,T3\W����k�/-����3�i~�bh�qf�~-�2�QI/���*��n%�����E�N��{|O>{Q�d��S�u�#cr�8V��	W�M��Xn;��מ�?~�Iq{Wv�ږ޴d %��_'5l��M�:Ԟ7�۝h䮧e�J.:z3B�B��͵P[��̿�;��ܰ{,�ѝ�]�5j�I�k�lO�Ω���&��>��c��-�����f�lP��[3�(�g��adHǵ�h�SZ�ld��L6�%�H)���!E�ʊ���vվ���������<�7�U��47\����ʈ"/��}`i��@���?��]�a���>'~�h��=C��0/z>��4PR��&=��{s9Tu�O�	B�uc�C�d�۽0^�����h��6+���I���NB$q\�Y�+��d��1�w:����̥�ĘD��|��L��"urH��M��,��o����T���GJ��}D��Qȡ��Ѝ|�0CZ\�	_a���6/1�;����Kq�����>3y/�l���~��迾��s�1k����S���������&�|�I�֔�QKI�u�#}rpSqw:��^HX����L��咷<^���nd��(��\J`�[i���J�P��h�c�s.h��_�=�F�`A��/������Q�]�6� [J�չPg^�u�jj��uW��~0s�s+LJZ:�P����2G�T�����q����l6��j?t
^_�`b�.t���z��q��䲟^�,8,i�(p9�� �hK'��^�_��+�>1��+�V�q ��G$�a�A7�����:F��N"�}`l���Ԇ<v�_(��Nޗܘ�~=�tz�����,�CM���(� 5@X�Q�H=p�^´�X��H,�R��Kژd��&��󿴾_�,6	��&W�Հ��}�6���\��<j3RR~�����p���T�N�
9)�s�PW�M�ђ�g�v��Ipg�v�2�a�� �x F���N�����iZ����l��gqg6�����f�7�z�9��Sڷ�~59y���i��P���Wv�0M 4!O
�ղ�0�a��2]� �b�>_�x2kd�����M���d�����i!WK^T�9. (�����rKX
v%(..���|��{W�����R"g��5��o�>�@�2U�T�2����=26+\�� V��5y_�͒��(4��+��fHi��fe3�Z�����kp�$���!��_EH �Or�"���Ur�
�fG~\�k�Q�S��Y�Ogu�V�at
�Ȝ'1�L��|�o���l�Q"����"��t-΁���c��y2�Gٲ�H�	q�������z�݄O�W?n�2~�et�{(E'+��/�J�X)Gz>�l>�OŞ���<��P������>	�W�B�UR�^W�ַ��s�YW�,[����2Wr�GZ%�ʁ)��q*�b��w�R��JO��p��)>�@� W�����5�ｄ:ƴy�>���2B��<޳'ï��s����ڻ��pʬ�A��o��u�'�p���=��?�J�
2��ԏ��vQ1#hx���ܨ�dL��h��b�>4�%����J�a3�o�Ƙ����W4��p�M�-����x qק���"XeN�
5�Y�j����׆4(�aO�z�~�рJk2r��PB�x���Q��8p�ٽ�4��^���<�n�n�I	^Ғ�5��S�̸k�����O�x?��0W���C%�7EB,���d/���6*99�飉t��)�k�pη�Gc��5�:�'{̓t:Y�7�1a�03�����/:b3?�G��<A�A.~�"E�F�{�i�Ygq��ͤAމ�ȇ-)p¬V���C��y�x|S���F�������*���;�ȟe7�Z'C���o��o����]Yl1<���8�i��U��"^�:���fw��9h?`i�9�����#ū��(��鐐w��0��t�|DO�u(��n��R�o�g�㍮	^�:f�ͳ֩��b���a�8��w΍B�����~������'9:G�����g�ѽ*`���g# ���~$�GwE���'j�����+�笡�=�g,>Oc"B(�>q�jD7��Դ�.Jꧼ�`{iUΉyJ19�bB�{��?�Pr�1�<�=�2�1���p��U�P�d����C�C�uo��zl���	#�������s<n�sO������>J0�1|/��Il���1�_���T��L*�a�$��Ye;�����u����k�p�eb%7��n�ޟ�o��|�$��"�&5Uۣ�?�IH���'��ք�äYB����~R5�������Տ>�ߊ�T"zsO>�r?��M��l�>|7��E\�O\@�h�Ό��aH��ڧ��$��D5(�/G)t���/�˵�ʣ1`��b�Q=7%XP�*{�!�͚~~ =d4���Q�]f׽FV���ѩ�co�����\��E@��f���<�nu�+T�_CͮU�� ~������B���\"$۳�\�{lUj�\zrxPL,h���s%�غ��f�TC�
$�H��O�^m�������Qa���Àa�}�t� q��&r+^)�dT�$���n���D#o'm=�"���������#�_v��[�ִ���w�ʡ�WF��������2A���m�]����z3�� �0%.����B+09���9�ɂ۸��#��s�&�F�)"<֐'���B�l�a�F�o��m�����w�ߴ#b��S=vJ�75���\��ӯ�yW�1A�9@�
�J�z�7��䅑aÈ	�a6W�	�M�.�ߚ8<��t�\SD����W�;8����-��D/���`��k4����Ž�������c��mv��B�����5uN ��� @�(w���twK�`yRT�!�~d�@���[��9�y��"�@Z:�U����]�s�^�a�MZۓ,��Xi4�%�.�D��HNi�vm��xo[��q�{��n���Nw��%�5eҿ��d��a>��8Z4iU7o{q�E�̈́c����>���JF���;��mқ���rل����-/�����zq��i�����v�6�yD�c�V���n'��@|�
�%��/���e���8��S�$���k���o��D�.�W	"������tK?�����iG��a�>�8���i����J�����%m�����p�!���j�=����� �C6�T�do$��x*m��(�6��>Ey�B��v��umAd��	�j�y�Ê�l�65�a���4�T�lYq�MKo���e�6F���эI	�=lf�D��Єl�.�� u�о�
���e��"��;�:S�(�j�^�!ơ�^�<���2���=I��A~�_�u�|����O��"��M)PA&8����+�:Tk�𔞣(=�i�*�ű��$�pRd�ƈF3H�t�Ɲ~�lC"����M?�/c�@���G�ڲ���b����*\��	w�h��l��7��2�����on l�fG8��C�A'���'�,��2\r3 ��z�V���Σ���44���ZF� ~�$Ӷc<z�H�" :)����L׏�c��˛��]�;%�c�Cj��&����1����n
��b�"����a�e-�s������� ʡ�EnMw�u��~.ρ)����Q���3��h��A�a(i���7q �EVa>@71�}׃�yV�!������ȁ>���;L�����^�Q��'���u�d9auU���[S�jB�4w'���V�JDm���BI�"oc����Lx�?6�n �
�:ag�s��~xH�<%���eOz� M$0~~�R~[9��C���t�"��Z9��i[K6��I�#��F2	͉�� /M��h��kT%�51�B�+J�T�������Д�-�8w�x�K����'Ǟ�<涠<?N��H����� ;c�/����֫���S�T}�\���Vg))z�p��HG��@B'��a��po���`��O�\��dKj�2W-j��j���w�ܡ|��$��UEЂF�^ n_�wTOW@4H577���Q�HR5Caf,����\����f�%����'T��f��q�	��0H�rZm�Φ��0�p��v�F�H�uȜ��G�A����p�sr�� :�U�^���t�
��`dG�=˅���:�*~^�2�,����b�Z��ᄂ�Ȣ�mYh�W���vNfQ�9R4��=�s+"w1CDe6F}JCՃ$��=���2K�F�
8����f4�Q�jU����]�w*2ɫ� t�9]�*�A/ ߩ�Zu��zE`�9B������K����iG}b8�5��B��r�w]��y�ht����W�<nT�l �H�2�}�9w�J�s�ڞ�c�JF����j�U��T���J�2H>;���E��N6c)?�
�Մv����N|Z�+���㨝˔|�8O�6#�Od}2�mhΌ�3 9Zμ�s�7u�	^ў�cF�f]��.	���۷�z�:N���b�;��|L�Np_�j!�`V����!h�u+8�>Z���Wyũ���9&�]yK�r����|�y�NOD䴥���z���m���.)��G>�S��x�Q�ADI0�]�]�����6�h�pShu��[T�d�'���gv�j^�Q�\�N]~����/Fs#�����c)��$�iY��i���R���u2�%X�іyd��)Ց�D"|��}W��?�PҮfV�o�G�7��=O�ߙ,FF��n�������̓�!k�x�F:[�����uȤI��|緡MK�f��+>��Jڤ@>�R��r���O����~��@�j��)K�e>��˼z��d܆�֫D4�#v�#��S�vC�fW�sk����hm9S/�_�
�a��+ �o�6W��v�eڵ�v0R�X�|�	�yϕ����f%�4� ��8�j��r�mL�uՄ|��#��Z�����Ð��}e\l�ylU���\5�N��͹��0>��t^��U"�[�L�uW�,H�����+��_�	`W���I�N%�_��aqc��S�3������IT���Hڱ��J�gN׃:�1��ca�7c��pM��5I<��> �������f� ���K$?s�'(�a����q^g�@dت3�fB�mnElr*�^���jq���R������*Ou���$�f�]5��X����O.�_h�)<?G�dA\-�
-Y��S��!<n��Q0o�G��=�}Y�he�އ8��+T�J�;��i_�:��xǎ���y��j7��G_B�$���&��2A���5S2�s�ʋk���wd�&"[���&�~zLmPAa�wc}���9l���I�c�	� ��eIH�fX/�p��n>���P
��v�v��֝LN�>;�}d]�c��b�����(�;غ�>͆�B�+�k�뫵�8�l��*�1O�s�/����c��a2�+e���{�,��5�U��Bl.[���S�Yհ�\a�vl�	$�*����?T�]яsz�{�(�9�ן�TL������`ə�Lb��\3�y�xj}�U�cZy�0פ�R���	�~c2��y��Ah����{�u�AXc��	{}5�����R��$���^��r�&��6��+�t��W�w�l�Lc�;�⻟���|����Fڦv�07:�����A��߄���2LV�e�P���Om���YT��Oܡ�>�(:	��������_ꜷ�+b��1�Cm{Zƨq��(����@�[FI���M�,IҚ��K�+�D�,����.��^u��:����^9��:pl�L� D��ntgQ���^.�8ĥ�q>�e�}Y��"��A5�c�,�A��l���(�R�y��5�_6[�*���|wrG�~�4���>y�o؛�B�m��k�#�Ph�f�	��3���Zq!�S7c�!JY�g��e�S�"ܤ�;�O���Y����gw�����ѧ���v��ms�&#��c*�b��3��X��|2K=���:��Y��b⁍����r�(k���+��9��p������h��+cyKU�E0�� {��q�ƒ�/	�aL=1���9����j���%��D��.X��p���l�̉q��ӸM�/�8�J@n>�1��.����n��v��6�8 u�۟V���kFf�RK���q���Qn�j��s{���$M`����P'.җ"��w�y�|3p�G�s�$;D��Φ�R"&�l�sm��ګ�1V�.�D�&�N&����<|��m+���|�RF¤�{&��?�j�j�����h���6���WI��;V+P^F���kQ��A��X��wS������f�7���"���]<�?��Hy��?�a;k��&����կ�@ˠ�q*/cԅ,�#[^"FG�PcöRCc[��J�z�ֺd4�'�y�z%D�ݠ�?4�$�{���}����^n�R���݉��7�T�4pR���
->��xpVڂ��J[\�_��m<e*r��!��?� ۺ)V��8>[6���t��Č�O�Z������߁vQ��`�SYXo0_��0��^|S�r�r�#{х�"��M�3BG�"����߃:?VG�Vn���-�Q��1�'͸��R�����`���4sd�É�O(��Ö����s��7`O2U��)����ʩA`Х��~{$��J�L���,o� �3l�p	`�Ȕ�����,S�υ=)� �Oe?�uI��l�wu7=V�X��Xҹ聘�-d�W��h� }��,���b�$űF��L�Kd]b�X����{?�����X"�@dx�9��v�����@��T
��hNL�+�Z�{ �΁�x��r��`:g��/ ��A��:V4��gB��
��ZJ�Z�R�׏��R����)���l���/T|��r��29�D�ђ/_��q� ��x
	����I��E�ڜ�.�D�Bߝ�����?J��:��]Ԍԕu�Bke�)?�4*j PW.��R����Rd����n�����+��'=���~����zju���;'L�]U}SWθ�?x����.q�G}���K���s�ʪ呚����f�*-�M��agVAKA��ߊ7��Nf�+g��ߗ:i������*�3X�A9#�%k^�h�_�V8��E�H�H/��3l��9�9�9I�:�eK�ؗ�2F�T<���?��B���9zө]�
mm%9K5 �4�5�+Fa+����8�V[�-@��bJ�����	I���\�lV��E)������z�K��^o�t��-��n�\��u������/z_%�P2�n���e�V�M�o�J9�aX��S�R��{y�QVZBT���K|�����#��e|��i�c�Է�NZP]�H0Q8�P����oC�ܤ�H��l�I\�R*t�
܅� 0����#$�Tȏk��m�ld�T@��$�h�13r3ɫQm����+D*�K9���=������^�(��=�hQW�6w,c��Y��092�W��r|	|Q����g	LӼL/<4C��m1ݱRD�Ζ��}؞$�љ~�<�W��v�z�p�~���K�%˕�ħԓtr���fL�ҝ��=���Lˀ����+���4yD�,3��h�s�~��_7U�;�ӑ�|��9{!	O���e�0�Z�Q�g!�b��c���G:�zu!�fvv=��K�r�R��15k��i/��+�6C��X$�@䯉�n*
���Tt4��^^��p��������#�����xk'��ӫ�X@�n\s�q�1�8#gԠy������IE����D�2�5�&S"�8�kxb������
�\d��/�#޺d�&
1�Ƿ:@煯߁i��3�i���M6�ڈ�,.�9\zN���9�#g�u�%�`6��(��i 5���γ0�Kv���:���P�X��ߑ���d��%��jnoɲ
�L!��<E��{�S]�I[2��b1�KśV���Q����qS��Js�@�u���d+���QY�id��5j��5oz�����.�c�aI��_�	^��_�A*��R�CIS%��j�c�;j����o�VKE1]\[�J�]��	��"�N>DYe�=Np�HwGТ�Ca����/�+�k��]�<-�`dFZTG�h��� �y�oZy��x��·�e���h���(W���=ن��Y���xq}SpP-;1A�4�� ȡ(����rʺ�,�@G�(�d�F:؉�y�=�i7�H���[�Bܥ�U,�(��SiD7�lw��j6��<�λ��߫L��:�i�b�kc�V.p�a� �~Ќ�T���>��+4�t�O�+���;z���ST0�� �Z�W2��W8.ܕR�B�e!��C��;��*_���h![���Uj:��u���Bg�f�0�]�Z���+�^�|���AKۙL��A97��v��(Lt��H���=Ga��h�d1�5P�F��c{FLOe�Y�]�m׍�v챮̏8�<�<�eG����ͺ�А5.4i~0������=q�CM7ژ�������׷I.��Dެx�\�����=��'
��ò��&9�1���j�+�vPI!�\���<;�
>�9�LҢDBdwh�50��T �~�H��s��րq��t�E���WUi]������j��xΡ[O!�i-*W���z�N��F:P�����|8�_�������5L�s�JB:�c$�UF��0[��E>��� 2�0���sGo�:��1A�k�%�|�K�
�F��.,�d�n4j�^Kx���׋�3�RC��� ڽ������!��'��T�T����$�:N��K�Ck_�,��+�eD�<BMCn]3�]G�9����Hf��^i��������s����?5�����L֩v���z��v��>�M�Q�4���꣤�	���h鲀�F�H&�Y��� ��Ip31Ⓗc�yN
��/YP����cؽMU���Fa\e����; ��N�Z�?����SJG��'���!°�>�k��%D �mraf��?���Ư|o'��I!8V���,!�e�4g�L�'�m�S-JN3P[ �D�p��c�ɼ˰�a0.�
��Zl�~!�"���LpKa��T�R0����^r�>F���MzJ�_p��J[xCغa��]����.R�s��Ke��7RI�(�d���8X\��Yj�"Y�.S�x<v�㿑}�J��,��mǨ���V�mQ�)2D��|>9U�F����Bʣ�A�Z�x��h	���e#e㦫�o�:�_?���e~SV_J��������v�_o��K�8Cxz���Bh��4(+�N,��t����=��e��G�2��m�@���5�r
B�ʄ��ہ@��i5�.�}.J�x<���{���f���+*6e�]R��\��0��g5-�9S�C�@�n����/� =:�;�>�$k*SM���p�!2�zC��9���e۝.�!i�kܬ(���T�M ��M@.�d9����>��i�V3j��1��>��<.���-<J�x���Gw���G(%��?���N 3�*ᩙ����� b�q|ԮkL��������/Ȳ�(F��KO�k�L����0�M���K��h(�J���D�V)7�kX0��#�M�1̒�-dJ�^%�GA��aoa�����W_���Nl�CQ�Q9N��cT��{Q]+g�p�5�lw#'�Gj(�
�y�'4Yp����1���V0	vB�?��Z�bI�����-���"��2{F�}�*�A�ąW��r����q�
��8�'�9@�-.�F�, ����Sy�m�y5��)���x�p�.^+��ATKH�+�1<8)s�~��m��L��`n��PW[��`��D=�>�V��\{_�Z���L�tsT��=�3x$��B��.m�
AP�~2w����m}�@�X��/6���L&�GF?vk�8¤�E�.,���y ׮nR@�heߢ�}�Z:����d!k�T
���I���HD	"���(�u�q9��N2[�6�O���lrb�0�<���Z>��(�3A�C�HW�-76��⩾�}��(��=)r�*��?7vj� RL9X�E� V��cgk�*��Xx|(��c{A�#��I��e��G#~&�Sҡn߃��a62ڞ���� Uy��)=����ѝHJ��|�����ii�uNMr�H��A�~�'�!��!I��Ζ���� x���;�s��"��Wc�X�{B"�N��23ԩ����EN8g��W��iX�*um^�������O�/U�)+���]F�"Ʈ�K����i�??k@EpL	��q��ǣ�pc76Ȯˑgd��w�/��\.epk� L��$ʚAY2DڼK�(y���3E��ߋ�m�܈1N��&����I}J<O��G>!��^(Vp��nW��Ѡ>�%u��R�{)A���t�O@cBP�'�Vq뾵BUJ�S�{~�!S���%{���ܾ�+|H}H'�J���J\3���!zJ�?����5����9��U�gHEɳ"p��\�������rJ���w>��hb�LDnh�T1x��j�f+�/H=ǁq�Ҷ �i����x��l�+Ll���3S��X%b�wKp#7_���V��4^/�ak��G̥w��-��F'��B�e������瓽�����!�J���q�qP��w�T:L�gt��3ì"�`�;�ێ�z��Y6��#�o�êu���n>f]�gϗ<�-p�Q]�P6Y�z	H��^�� �9�Mb:�m���*�O���r�~�o��v�
�lgg�0��q逡W���~�0c�������N�A󖋠v��+J�s"�s`��� ��@��k���٥����f~�TO|��G�� �;ַ��R���	r�˺$��kHQ`�9�稽�D��rLJ^��%���V�78|
�������+K�Hx�<wpJx�	�Źn ��� o���h���[E#��di)a�N��lY�%S������Oʟ`�.����Y 8�L��Mz�)c�ǉY���ӈ�\Y���ȩ���h2�ܵK"�[�v��)A�����"x���b>w��Nj*7�YV|S�3x.0�za���ጠ� {�B�[�-흗k���Y�P�C�(����x�B�'�/NQ��*"@��M �-7lǘ�nAD{��m�I׿{&.g�J����{[�����z�&]p�<Dе~E}[��g2��W��7���u��C։��jM=^1v���:�81���k&E�>b�'����iҐJ�ڿ�*��G����Ƿ�|�d������42�c�������@����J���d���5 
�����"����2Z-�T�%�`�d����2��mj��ˋ���K�$�o���F����	l�,���'�:V9b����%ej����
U.W��O��R	u�Ow����!*he��Xی-�Er���V���R����O�Np�/����h`�vD�4�u`EGK���a�8+���`C	�b{�=5�8��IB�ٜ�$#�X��'Y�(��0/��7ŋ�3�0�F���)@�<���$���8�E�r��RE���|3H���-���1�r~��	ƝO^eXA1��[㰰D�ݝ�a�ML�������@$4��Ix$���8�¸1�IJ�l�$�T?����*3�h��fXI��V�d8�Ħ鰨/��Ү��}]�'[�l�h{yUdZ@2�7�Q�b�k��i�X�J)�nc���(��mb>x�}��ch�����8P�I㯀�>hz"��rE��٭��>ñ=�D�]8D��!�O�ߤ ž��a�/��Ģ�?�8�)\��z
��>w�9EX_s:��5sm�����l#��U;})8_*�Kf���t�VJ��`��k+p�k���Kvn��M<���!���7,�l;�r�U{�]�̿<K���
���W%���Do���7�3"i?��^���_y�J2nCE��n4�*�vq��A�~��fn�ac=�߆�5���^�,�܉l �P\֍��J�t�&�>�9��7�b)���YrCl���A�ծa����#�ˮx��9�c3,�kf�9ܖ�&s0�q���l!�=�d�Le�����b��e{hD��h$Un�:�b^G�R�:20�m-�[ö0VM�I˄��ĸ�z��������(PN�R�h��#ٕ�t �E�|��;�W��영������d��+��٦Ԅ���-oEh�c�K�Fb�0b�eq�T�z�2���,"?FeTO��v֫69��s���\K/+���у`����8��B���Hd����2�ܮ�b�<���AwwpSΖOi�[9}ڞ�+���#��>��)6[C{�i҆-RR��im* ��k��g��~6�6Eh[�1��,x�6��L������Z���$��q�ˊ"���5��L��N��N����j沣O4�`Oܟ
���| �/2մt��-e39�ݾ�uo[��n�R��]�_�1&=�����h�[_V�:�-�m"��gU��`��G�2j@\&��'^j�`�y<�_M}	9]�v9� �;/V�h���>g��D�.�����L��,�."ș�ľ�x��ʅ��˳GV�a1a�}0����횋rMc|E���=�Jt�[U�r�(ח�&�m��Z*�g#p���'JY�7�H͛�7�1�<���$I������+u;�V�0o`�-#ƳqJ�/k��W�{����L�������X��:�6��ka�bw��#&��XZ��N;�S�eoV 5��{�P�ܾ�AMgD�j���9��Z߅2����ޣl�����Q{9 �[�<�ۏ����&J��/�jכB��;�ސ���Sq
�Q�əǡ6��/�n���;�Ѝ~�O���MX�*��%��+��s�nˀ%$��b�`�݃��H1�J�A�:�Z���'�h�	�
�G�ه�P>)��|�*R��N�Ї�|TP��_c�K��C��R�˛��ʜN�k���n[�D	�EC��4f~����a��a��gc[�D��uD8�^"�!�*V�]�w[r�m��:T��:����G���[�� \:n	��`���Ey$���O���ީ���KO/�X�:�F�-���7%�I'Ab����߉ϩ�D A �j,;�Ŕ�tL�t�:����*���k�.�ӯ�(��]���>�T�:�g@��H�wJО��AK�r�6,Ĳ0�/��6h̏�����B���i�}e{Fyd�'@�&+o�,$����.t-ޅVFL�Ր:S&�4 qu�����̵쩾�Z,���H1�፥p�!�0��˴���^d�4k��GDN(�\x�}�J�����}���� A���_~Ƭ��q�T�2ꅀ�����^���P�Q��c��ʷ��yI��y��A4ﺎﳐܴ&~ĺ�aLXx�,�#����j��y�/��/A<�\G���L!D���۠S��8S�K�B��~��4���}?Nh#<dv;�Y�ܙ������Q��I��m<��ul���?�$��+K>"�_H)3���G%OT��Y���̚+ea��H�_u�|.0A����`(����D@�0l��g�Ĩ�^���1�!��U����E�+_��!͆��͢#̊d����]��E�O�G)i�`0�?5����Gn/�(l��|�gv���
s)	�}U��(�����DŦ�'^;K�9g���]��IİU<?D�.|Dy�d�Z�?n��/�,sX"*C�����52C��2?�j�a����K����|� ��ڽ_��n�G;�����E�>Lݍ"����*E�}_�<�����`�+Ch����P�Mǐ*���^���a<(��Tē	���5𒚆y�Sz�0��y��s��O��:o��y������@�A�G��{;�i���5\`�	
���&ר�`[}�8<O�nV�u��؄�B�S��HM���������g� �����Pc�d��	YLf9HLy�vp��J�q\�eV5�S��d�Ky�y�A3v�U�m)!J	�󴝩�~�4��l��A����+�ɪ�bT���Sĝe�A�r,0����{�݆ ��y��aD=��[;o=����@�џH�T ��B��O�}���- �`�	j`��a�ik&�L�Br|��{���.��ªѱ���f�FR���
X�������s�O���-r��������NO>}f�F��es՗�g7)@>��1�������_�����@6�v����A�7DXT�*b�c��W2.���,�#�֒�Z0k_�*cp�3
�0>t!��@��:LH�
/���3��`m��D���{"�안{7b�m_ā:�*_�\�\��7� �4UU�R�c�AaO����9��0�u���]��օK�~�Z��&1�S��v17�ee���}��rA��GݾH��,���	�� )lU387�f�@w����@|_��ݒ�{%�'�O�T��A����W���c�ZAUgr�R��#pr�^%|�*5<�n�]Y���;bR��BS�q1��ۍ�C�k�o���B�X��3��>y3�ј���Y	1��+M1��4���gOH� ,������K0���K,x1t4H
y��ol?̦�[��i ;����?F����K�x�X�K��_�����#�a���
Q��FV��t+���Ԧx���/���� c���z;�{����g���Q���@�
���R�O ��㉞FjD�G-~��#��@��o_eev�Q�+�6ޱ�(
������c1�.jK��wi���;×�1fIDf�)EJy䶭������fZ��g����cjyY�AF.�ҩ6��/ ��X��Ob<K"O����x�gp]} �%4�ŌG�.�4�_2���ٔ�c�Hf�!V���ܞ?P��?\����-m>G�4�2��2
��eLӃ�vfߔ��� "İ)�5�d+D��;F&NRK�=�qH$�s���-��Ժ�1ˣ!��&z���1C�S�ɵ])�Z�M#����t�f�9j�^J��� ��O�m��<�I/�JАK�#Ul�H{�pAw��qR��R�P�m"���+E5h�,��ǎ�K�?�N�+D�.2�_b��#��
þ�bG�����8��26\K�u�:I�YX������k�n���w��5�����D���uCay��7��UFctr���=0/4�,�퓦5S��w�t'�*z��$)dk�8/r�M�Z�({M���.B�[t�����9���mY��NU���G�"W��B���>��ZR����R�W�[ �	,;Ռ<��	�	�;@	=�9�z�oS�lpv �8"��4��=3��F�-�	λ�(����4��?0�
砒͓���8}#D��۞�&;���л�g�ӏ���c!ctEwZ?q@a{����Pu7Uގ����,�{9��~4BLlxs��i���>(C �f��Z|uZ���k�qY������ǿ�6�0I���n�������}�XY��AH-�:�Ka�������rg\�K�Q���Z�O1*RL�b�v\�~E�H��ۀ{Sy�N!y����ύ%���dи�żP"�����v�r�#f<����4�S7�����e�/vy��@U���hӌ�m:rcisrDz�Pz�ٮ7�U\	�v����P
��睮u���&iW�Õ�n�T��ۭ  ��;�������)�1��%;����l����.U+��f 'ܾYX7�Wn��$y}�ϡ{Y7�Z�96aд�`�5V�tk�}q�Rr��IaY�+�ʏ,Y��,��������(�F���5T�m�(R�>)�ę��V�?2�9�F
1�q��m�G����~���"U6�&ΗCy��3�b$?��u�z��L�\��%��֭6̸k��*U4�`_�WsqP�D
�	|E�
���ͻ<� Wٰ����xp���[X���c��hÕ}�u�p��c� �+͑��ʪ��4Tz�'�>t>�O�z���}6��ЩZM�J.��y�A���2rn/�!-��`�Γ5��|�p*��~ �Ȇ_���|��`��t�ڦ��u��I��\�r���򪪷T�=��~���EȒ�i����mM����������}P��UԘ�7h�ź���F��W��0�%)����rc��-�/�v
c�����ķF[m�a�EJh���:�2��<�f����P�5�s�/:(���F����r�$����� 5B�w�C�γ�ǴuGS�eKO!HfBR(�ܮB\_J+:l�D�lD@��ˆ�тP��I��(�;���h�4D�T����!\z*���Sm�B'��1���D �Z����o��["����J��m�4���> Ij���Y�/��	aƧhe��7�%��<N�]З�Ě������4������y*�xj���^8��$�]�^ޔ��F)���r�o���w�)�8�(��\��&G�/Z@f�rCɘ%�Y�|�52�1z�A�����p�n'�W�2p@�Ϩ���v*)"Ȼz��a������,�Z����N�u�)��ZB�g�CC��)�v ����@Kx�B�N�O�p�8d�J����}~UW5UuriJ��/���j�ȡ[=�~�3S�햑z���sop���]!�*�G=Ÿb{I��],��.�N6�O�mѲ:�qk����T4�X�fZ���k_�����8 y	�'��}t
����z�w0��&�ea��xe}p7�`Ĵʗ?T���������I�B��)�\]Azĩ�C�K��&���	����:x.�6�z�Y�ٓn���ɒ�rī�7��܈�
�����u^�f��E�ʵ�%?���,���/� @hd*�>f��v�ZV�
��$��=�E)e�%��p@b�úZ'�o��>j�(KSD"��[{���t�`���T�Vg��T�Z-�Y���f�Vs���_���5a��6��F��kTL����x-\�o�/#�eZRPnu�%��=k`�0�XdN���ܺ����U���iS�)�/A��v������ڲ�ǁ-mY��p�ë�E,�~�U6��Q0����'/��7� R�'1����ap)�趗�.)b����I��VY$v�Y|���`��3�T�~4���D�y��$mY�i\oI�SJb��3-A��?SM�bj̼�\M>��4x��$���	a]}���<��\ݪ�r�M��U}C 5<ЫH��G��B������K����x��"*^�B0�KH�J�<@���cѰ�s�yB�Q��q����+�[ �&��K��43�H0��vػM[i<����j.e"��f�ɞ��M.���:^�z��V)bfN4脞
�B�lO���&@ s�m��w�`��70��4⼇��a��z��&����D6���؜
:s�Q�v�l��S�Z�u�b`A����չ[��|����Ԣ}��w�[�)���96/5	k�u������d:kg����;��4@{�Φ.��XP���"���6��ko˓A�s��K����8AI](_(�R�Q5�������G�	p4^���7 1��8/��i�~a��^�kp�"����}���g��C�ֻ��^�v��+�l8��t�$Hv��\@��L{W�Bv������]�9��~��V/I�
����a=U@y�a3�D�h,�7u����q�}���聮��ok�>��lP]�η��؁rY�՟inz�rT�F���O���C%'	�S��
)���j�2k���7C��x��m��/}}N^��c��Y������&Ύ���).���$V�%�ZJ`�j�^ٍX��=��K<������:� �+y ���qM�^k�`r��Yym�!4�/��kCR�-5U��"ܘw����I+v���ޜ�b��%kZ����>q�;�'R�`���	��Jdh.�8LA*.	/M!Ɍ�|�d�z�挢��y|�1c�v`f�J�Y��B��qj��X��K@C�W �f�D� }	�Hr��z_���Iv��T����q�$eR{f�g�hSe{Ki�ql�D�˄�@�_�zƮ�0��Aar�1U�(X������)�[�f��:=�&�X�_�CJa"��`��|I���34e�X���5��,u���I�a�?����k���<)�n���9k-����8�@��a�֎��)�4���ˮl�Xa�a�n�!t�ca�ī�Fӄn��%D������v\�K���gQk���Wb��TsuV��ό�'Xf-b��V�H{������A _;���#�]KI5�J�5n�mW|�����\R楚�S�M��c�E��BH9�Q��k���)q�o&:b��~�_�	�(�ǰ��i��No�w���?�,�)��G�[�C�] /q#��kñZR�D�D�@�T7boS�sz�<�CS~R�^r�*�o�U�xI,��4%Q�,f���<��er�ٓ�a�����5l���4�̂,�L -��>>�T7��AZ�A��B
�Hb���^��,�rZ0ދ����:u޾������V�K�L����A�T��ـ3/��b�ķ�
H��8�S�8%vaN��0�JEr�9�&C�h��&���ߐg\�t�E�m}�g����_���=����m�zɒ�4z�YZ�wc�h��}�G2SE��Lx[�����+/�H�s��=f���_q�MH*�w��\��7ESL��]�5��JXt���T;�d#�(& �}Џ���9b7ţqI868h��9�A����*½`���j�x�#H�����!�¦�T��0b\z��5�>oع°t��"%���P�*`��Y�m��@��B� �*� 3�t��1�t�e�(�f�'H4�V1Ah*���4�,���8��n�O��Ě$�u�K� ��3tV8_<rqO ��;!�g�ִbk�3�ˇ��S;Չ�{"$ܨf��S��܏Rd�)u�\��fn��K��"��d� t[���9����!8;��l�c�O
���=�巉�3�P����L��0m�`_��59չ�/�'�>��3rm�r�X+���+��j����~���\��kTrv�g��� �t�=�ύȼ�[����)w�MT���m??}%&��yA��8s6X�T\<W��~8_ѵB�f��΂d\�~�[i$�"�7�t��:3uV�=�ɸΊV������NA�Q���r[��Lm�`ՈtM���a~��*|�%~Җ��ʕ���(���¾Z K��:��7rz��ߦ$
ʠJ�ʪ�{��^��\F��;U�#\&K�'��Ҽ��ї�lƕ�wU�;������A��|�;�J��Ճ�t��l��#^A�
3a��lI��Zo�v0�"���H�J�@�Z�bh5J�c� ����	�a�?��}�����Gn�ܖ�ҧ�`*�����G��4�n��M��ۤV}.�g+#�39.�	�Xެfآ����^���s+�r9��I1Ӻ~��N�+S�w8���|�(�x�0]�W��|'}�[�3�v��	"���a~~�B)G�ț���d���+J L2����\s�;@�F��B��:&���$Ш��>��x$�Y��Z�u�Y,���&�Cj��bݕ��q(���ony��F�U��n�9I�f��4�9�����`j�.ӥ��Ut�jU��	c=_3����l)�ٔ�5W^�����ń���E�E:?�D�g�*�]L t˲�t{���g<	�2j�I�N�Q���"Ve��+\�R`ҕP��e�����͂��ô���?s!�R����=��5��ww��u�g�cU��(�B��X8��g��|��7&�>���Y5��������Q09.4�)�c{"@��K\��!D���o��L�a�u3lX��z�LٺL�W�-�.���Wj5�����V�X��r���?�G�ؒE�"]��RC7 Z�zh{��gf��&����o��� Ff��O(�<:�S���a��0#d��^G�˖����7��A��>��黋O�c�=���ʝ���[;pQV�MF�w�rG�&	yG��X���	6|��@��ӟ��)l�+�*|�]�~d���feu�f�l��x^eQ]��	�'U���������J����������8��6�9�QPB�~�r���>�K?X��x}�_!"�ǧ�s�]��������t�����. *��Ou�k������c �ZqS����
�1UU2��s�傓Ք��IScn��)c$z:��t.���1UjR?�vu�Ay4�!���P>\Ys���k��Q&'^��^OA���`�M��D�:,�?��u�t�P(�|���s�M��x4n"�TC�������@Y�������q�P�ib�v$a�v�p�ܨݍ����RȬڟ���>�l�{6�QxO����q���Pֻw�o�V��-�|h 7<��"l]��,9 7�P����^<8�P�1�����GyID8R�)���'�-�T	%��&(��u�j��N����� ����8�����+_	f�����[W�[��蛽�[���It'>����}�4�B��Gm�r~�(���>�V\���xY<� ��j�mT�шm^�e+�U]2�0_|œ�]�ݬ7���gZ���2�0bh6�uil��,{lpL�3EZ<���c������f��V#�([�	!v �� �e� ��dqCk��c��'��"�d o+%�a{Y'����f��l rJ��|,w�_�^����H�W�祼U��I�� #.�:N����d�j����c�"|���+(��󞲖3�'<�o&gK�wn<�������&=۰��~q 1��TG�|UΡŅD���5�
�,56
��`��	����,o�]��	���Ý��{ݐ,��<m�hWU�#��Z����s��	N�\�e�%/w�_�6�L.�7ȑ1�Δ�P���+��� zDN����,��R��/�� �0}0�i�
��r�Z#ڇjD��ޤ�3�c��W���E<��C�*�!�6�vĽ l�J��L�b�-�Q$z����gqqN��X��I�'T����j��֍-l�����[E˪U������ߨ���B��O�}p ����e�",0�}&EI�(��f�dJ�.��ҭ �����)[�����0�-���{5���b�A��f~�
8GE�d����� ���Hn12;�\X��Q-���7��I���(柷Hy�V��ܮ(��Y�:��n������Y5�tH�j�uiJ1�v_�P(��UU��:9��$l�D����=<֧rټ�+q��XŊ.X ���3,��![���2�Hr5ʐC�7+ٵ�L�Fԉ+PL�����!��>������ $K�t��1w��:Z���Ȧ�L�����z<���^/Ph��#O���N�7J!�u>��H�����[(%LgP���D4����CV�����]�����\��W�Q3R�(�i�
����Gq��J8�|}�MN��&t�����Y��P�𞿱�o1���蘬 /����U�5c��Q��<E{_@wv�#�#;���x(:@��.l�~�0���}�|M�-��l(y�h)YR8q���@W��K��Y�uM"�(9V))���ֱ��+ڬ��:�����-ƌz߁�"@'����RK����>�r<�3�r�o&��%,��EKas���Od~^��3`����!�g7 T��=ޕכ�\*�᫔/�H�H��r�j����f^�dV�/�[2:5bD�<2����^_� #ôx�j��_eǼU��%�á�o;%Mu ����qj���=�S�rQ�k<�+yFa1�K?�̦U�c<���ٛe��h�"���I�G�(�b���)���*�r=l��R� W��w��,Z,��H?.���F1*S�e�+�8��{�멅�����w<��(�ƥ/T�/�3�X���֥�lǿ�|gX!�e[�z��OA4�gi�S�|&PF����U�e���{�xF�X=A�b��`�ؖZs�{��g
|�#u���9��p�0`��"K�]���>����zU�+�lE��eZ<����sF�A�����j����د?7�σ�1o���'�$`���c�Ϊ��+��B��T�r� ! 4�{�AX��SfQ�z%�}�@�l���=��x%�?��8���
k��{��K�	����<�Z˓:�����'���'q�Ja:;����/��j����Sq:�2�5���r4_�����^1=�e���1��Pr՝W2��l�y��e,�R2	\:t��~ K���x���.�-�?�x �V��in��Gs4�Fe� ?�-��c02S���	M���B��$m&:���4������,����?���w�mNm����%|ܲ�n՝+�\6��]r�G��,s�%��+����A��y��OV�)����W� ��Rt�@�K�,�+K�@c�7��e�d��,�}GN�8�S>z5I�/j<"��~���H��R� F�,O�T�*�i���AD��O ��D?�=(MwGq���;�������8M�^w|"��\�x��y���1�-՟�v�"\��nb��t���J:�F"iKY�,c4&�w�&��X���,t��!Bo��^k��&&E�2�F���7-N8�[��AD��5�E���r��W9�{S��cI�s�I���7���6����21R��.}ҡ�K�P�A]W����LI�tJ*�XR>"��%zn��w��oPM�S�h=	Ɵ�C���Yv����So�se>>��y��k�d"�@����}����j��k���Sq**��>Qhz�ӵ�Q#`<�����\��Y���,��2 �b��LZ�� ��	0��|�X��eȻ7�g+YGM�E�S��v��
�ǜ�&XCʐ�kq�$���s{K��%����(��w엡��x>p��n�
��Ve�&�g����q����HIH�iQ��)�01�X���*��u�#�l��#3?�eX8�o�ŏxIc5q�#*A�{O�E��W�W�.��9:�p�evN,�����\_Mi�2�o�}:�ue���[���Z�TE�^��4PCi�8Ŋ���l��#��,��Z����:1cZ�N�D2u��������a GN������HFsja+�}@P3L%�Y���[0�h�MǾ���I�8Ҫ͚iJ�$2D�6���iX�]6�G�\�!��a�����/?��;�3^�Ki?�?t)+v{�3��&0O>M{Sc�5�U��H�[�'�f���z<��l��Q�>�5 ��ͪ8�U�Rz���Mq�
9�. ?"� yP���hIʱ���<�4��e�����|��0oW\��a�[���f�v�-%�n2fݓ��K��r��K�A���f��}��FV���^L�w�_f\$B�"悙om�N��}����H���/8Y�Y+u�QH[^p}\#	8�kd�W��3�<�,�#���R��
���ОT��>._�G/{`�c�O�� �P�{@��h��]!���;O1Q����O��m,-j�1��b�[J�.FO���%����cʛc�H*䒕�C��!8�6���ǽ��m-��0�%�̭jW&�E�5
��r]���\����$�*r��:N��Y��lъ�^�R�*�Ƙ����ܷB���Ƣ�&�OT����Ur!S��
�Y*S��xSO��ﰳ#~$�U�\=ğF�;ȃ�+�s�:��&�-�_��qn���h��H�V}�mM'a�>��~%��\>eQ�������V�;��%�n�Y�8_��yo�眆Hk�=Co �f� �ʅ��Fl���ueX51������Q��C7ưcr1�L�%v[��GY�9!WV�3-	=x����8�@�4�`nb�a�����i#iUۈT��ӱm?��p�	hP���|D�L���A��Q*	m��<u���vљ
���B5�7lKg��%��E�|`��)�¶}�6�O'��5 �\`��L ���.��s�łT��EE�@/�?ھ�],��D3-�'=��6px�A��Q�+I}@}��MTR�g�����E7�d�>v9�24��޺`ZlH�}��h"�x�d��X���h�Sm�A��$����N�[�b�5�����(�O���=����Vkȵ��K�AE�I��	��D�o7���$�Y��)/��p��i*��D��f1N�E���yGR�Y�+M��[S���ˀ����﷫w�8��ӯ�ڟLG#&�'��1",��K�}Ԏ�]�!u�ƴ*1*HU��NS	Ӧ[J]����w��ӛ��%Q ��$Pֹ:�.o5cT�+�`�Og���F ����˽%��~[F�
#<ugI��'.�؃EG���.�T`��D��a�\��3}�x�������قypy'l��rH��l�g�n'ʃ���s��������߀���5��e��pr��n�eDl��t����2'TQ�[�� r��m��nN����	���eӂ�7���}']c�{E=��i��Ҫ���2�jf&0�1��Ϣ[�"r/j�#'�b[�B*,�$T��|Bz�7��qk�V�D������Y���d,"W�y������L�)Q"!�O�)޳I{ju���%���܆��~{��F�R���$:�9�E�B*���2j�:�X(�뿹��S�@5�-x�^�QpcK*2 ���|�4��,�d��}�'�!��J�j6�R���4(4�M[��(��tt{7[*�M=]rf��M��gh-ga����IhUsT͟0i��k����3���
܄/[��x^`}*(��T��ԥ�3u4z]���jl�3����yK�<�"J���jA�����N�a톘U��؆Nc����MaDo�	�R��u)H��/*b� 9�tl�V��$y�� XvE9�f>�O��ݯ�zC�Қ�l��q�~}�4[�� Q��N�	K'
oB��VΘ9�@(�.TQ��H�y�9��N�M���%}b��4Ph;.��W>@2J��&��w�.~$U��\?�u��x�V�"$�O/��޹cE8M	��K�'��!��,-P<<�{�m�^��HNߦ?��wAC��/�>�G
�$���.p��T/($G�n<��-1�,;�ū��|��!��� ^�>������ �0����^�?����}����)�W�@��n���h��ᕹ[�+���-'?���%E�9�^�	�����Թy�D��=;`a��]y���g�����i�G��BY�1Sv����ц�L�ۭu��X��������YW��JBbiҪ�����C�~t���j�o�'|&��b�~���M?����{|Z3�sMA]���B/��eڿ���ƿN=l�7!�,{֐q�.��k��+����촚��fc��E�$	,���*	k������֓�GI|�^3����B��e�}_=�V���A/���u�[�(Ɍ<��6<��u�'�p|guFDH|����b`�}II*VF���RH���C�@	�#ޝ�6��Ⱥ�� ����<u�$�@ǂ»��d�Ð��<��<a�D�z����v���r%��NP�;����X���K`��/�r`�C����Lk�P�����`MQ�}��F���5�_�4�N�������ޟ򒮞�n�M~5�����7��|�ݾ��\]�sݼ�|"��(�_�Q���H��\(�y�-�N,g�1eC��"����1v�Xi ŗ�Ĳ9u^� h�����J��0�'���
Ԃ��O�zuWf�4Uk��x��=c� !�~�)��-�k�4��8��	�y=0ц*���Ptrj /���bQ>ǭ�
+a�@\~N�<��*��a�n�O���S�]��������f��ܻ�����J��ӝ(.]�>�ȷu���:�i'b��Lg[�����^��ܧM���C#l0gb�&m�z�-7:�E�)Xy��1�X�8��6��)���������'����Uč�^�j��E]���/�Тl�[�Z�i��� d}FS|>޶b(�m�C���L�>�jW���iy�j�|��]��<�5�҈{ 6�)��	�'�Op�sㆧ��i�]S�3�`Đi��P�!�⠏�j�DJ�TAt�;��6�g�{&4j�$�\k�O(��8S��'QϿ�wۮ3��������x�v
��GV=|C(�I�^�7@��VmU4�R�	�Me�13�@GM`hӄ�)�>�(H]�{vc����V�����8��k?a���щ:I�L�r�C���:s�{<�̜���lf�B�b7�����&�94jN���_��u"Ƙ���R�w�79���ƞ��A(�Y�8��i�h�B"u��K��N������V�~�DEm)�Gׁ=�P��
R���~���k�a�^p%8��ȉ<��<�u����R"����G���?�^�{��:��ma��>�48v��lZ]#���}Ok=�Y���i�i�
�w1���вh��⫭q�y;IP��{�m�������&]��z��<��Cb�-�8)V����5��ͧ�z2��VՀ�c��1o�fF��
����׈k3f�.�w(�mODa�s��6�����\��v���R�� ����7>�EAʭ�se�n�7�ޔ!}N�g&@�>%���7�C��#�S[OB��ۆy�m'����DS;�*���'��o����>�a��W	}j��(7�_`����M����{J��g=c�P4�3��&�{ؤ}q�ҍ҇`�ã�H���tuR�\ۛF���F���U# D�7ۮ�j��x.o嬡1���I�'ոp�2�~c�[������5HPbq��g�;�y�� ����5�`5��ΌhE��i��ݝ�7���`��v��	�$|*.����(��ET��x@gb=���sj_'��*���M;�&L8oнD$�9g���C	�^�WW/ꅧ��s�Di�aݾ���q�8����+9�k��
-�M�j]|�<�k�������U��rj�_�9�i��:&Y�|ӐV�0PN�*5���r
�� �u��f�Ѣ�xY�Tq�P��BвKPH�x����d����Hm��!���o��K��,+!#�~��3�IGE�<5a��iggyļ ��BY7��T�i}��a �������P�:���R2Q���`b��CNw��	��3��ИէId����zj������o�Hy��3y5(,�K7�ʎk�gw�;����y�ˉ�!�
�4�/�WH�/�0c�U$�|�P˻��gvh�����]��Ē��M\����FC�:'�+G�X�Aq�L2>H�Pd�'U�m�K21��
�{zs�:�=��rq?��t�G�'���A����<EA��A�=�����.�
yy���%,%9]�=:w��)�	�b��r6F�q��R��.���$S���%�1v��b��Ƅ>�n�[7���h�s�dʊ��&	�"�&|z8�ܣS8�����{�m�5��~OC���I����T6}��f��>��4{X-�l��{!�h?�w'r������
��.�D>����f>kJJ�ы���;�~�8��]}c�(��i�)�?���;ơoO/�V̒�����J��L4w�5�ؔy�P�8	�x�g��7+�8�G: ���d���Vf���0��UЈ�\�҅�~�'M�j_��QlA=�6Y�U�x���D��SyvW�j�A�x:�	=S��)	�!ӞmGb	W�4�G�*��lܼ�U���x=���o�9§b٠+��#��&�F�aUND�d��Yr�g]��@���Y/�,���8;u� ���7���_��4�pYڳfq� ��N��|P!Jd|����X'9�Z�!'�������%������gz��9���I�*w^�yv���L���L<��1L-q�R�Q�?\Κ:�Q ��GS���Q��YI��{��NZ8Mc��&���k�5v�_Y��A��kd���ʥ�f0�l�пC٨��9����{.(t�5Y���'At��]L��q ��6A�bQC��k�g YL���^��$���p�#q��9�~=X;�x�|��1�D��zC� P��ٱ��	;z�c,����H��WFbEw��^lG�`�xZ��Y��������<���_���ȵ�N�����yY�����VA.u��M-�Nq�{)�7�AY6�CG�V�U�ɴ�Y�`C��⺷I���߻�4�ؓ�T�$�2(���S*g$�>� i�*�0g��@��޼) ,�J�+q:����w7��_�h��W�WZ��p�J����	�A� ���dٶ{pГ��cH��%Ϳ����^�'������"���!�-.����7�56E't��M֚`r��C*��h�ծ�U�z��O.�p^wE�U�ߥ�45����)~]�y���ʨ�-'�x���|���T�r��ns>_�񐆑�;��?�m9�}�c�f�$_G�*���V��)fȎ8����cbs�)H��W��i��r�މ���Q�q�S����+��o�����c*���\�]!�x�q���9G)?�`+��$L��8��X��%�v�;��>57����T�$�2�ݡ9C��3-�u=�P,Bl��s�to�W��p������rF����M�π�0��}t3vTn5X;�B<�lR�V,���6I�\Hq�F;�P��fZ��gS��`ң~��m�~A�$'�Y\C#��J�ꆤy#�yx2L��|�Q�
�h�cH`R�2P�<w�.��&H7�����@8���X�1���t���:�| � 7Y`;�2jG*B|���	E�L�4���f��v�I.Z�8J'��L%"�p�Y�$L�ճ`���;�`Kk�``����A�<X��9�$"�eE��셆�r<�kȧ����c;л��B
�n��Lb�c5�Ru,����6>�|Uzz���;���u�,{�5x`9Ǜ��,���]�_u&GX �Ȋ�œO����聻�f2�/bϿi-y��:J����io�m��X{���c-���;gW��+JcpƹG���o��;�9}��x�4j�.�ƒ����+!�ڴ�{�E�_��UbI�b����ϩ��uSD�n�Co5�/bJwq	��xֿbG��t�����$�s���.̊?�1{��ר'�^o�r��#� l�z{���Y�-����;p���wGu���z�Q��`��<&�u�_m�X��5Adש\���A�\ϳM9���|G�Ι���E�ο0�\Ϛg��
�(PQ�hJ� �O�eV������u�eS�b�25��!V��,!a�p��
�	�1�G��#[��-_]+'c=��i#S�/�/���oX0 ز|�ީM�~C,��������z���u��߳�.J���a���*��Չʹ��?N���/:X�@i �\Ii�ݩ[Lz�aI���G>tW���y��v����"���V7���5(�
���MC4�)��r��T\��nL��4�>e<&��~��p�ߴ�j:l�Lq�ys)�w�z���{��J]*��S�H���=+xN�m�����؋NY�J��neuBw��eo�fY�J/]N^-G�0�����8ʽ�7b�u�x}��C�b��X�p�I��h{�uIH����E�=�Uq��q��=��r��Ͱ*/��?Q�x�+�}(l�o#9Q��_�(\�+������|���x����`a�I��2��D������簨��>z�.��~W�&B01qS�FU��$�(��r���nd+���� |Bɥ�1�#C5�&
X���!�-�ힶ�S.bk�<��S�vO��'R�d���r¢��#r�ENB�}|����tBm���'Z����rݴ��?��i�@��3���Y<�a�*�v��eٔw �V�k�@&��� �P0~�8�65�@�Mpj��ws�-�Z���	ʻ:~ީ��or3Y�P���C���,h��(�>����V����{�����o���%� n�2*q%î4�2�j(�Z��l�!JLS��c�C��Eqjn~È("d�����3��9��2��q�|Y�$�����q.�z0VD��:F7�����X��1����m�d� � ��3�c	9W��۝A¶��L�8y#WrRæ��p�*�`���eY�g�vrJ�Tk��7�cBm�b`	���$~��:�N21�jǰ׎7�3��N�ƞ��Ȳ=@���Zhޘ�?�yFL$��>�|�,"��7ڇ$?~��Zu��dl�f�_�~��2!|���H��2��g���y_=jp��ߧ��4OE�J���+\�66�R��%p}��$)�Lx�+��
�z�ރ����I�dsh�A�h��~�����"I�a���O Ş��|B��ا�U8�UA��.1=r!�?��YuKx��j�Μ���n娝	��8#ͣ0�[���FX��X�IA�8���#ީ��²��ٞ�^c�Ц�
�qO��]�ԌLܹ�� nl��ޡ�g�6��˗^��nᅷs9d{|�X[�x�Ӹ�Cn%�� �hz��	�Ǡi�Ի�ӎ�h_�� ��=��K�3D����w5#�,ڷ���9�����2j�̩�Q��	��g޾�S$���C8S��Y]9:�魠�����$�iJ�����EE�bZ���nG������m���m5�,V��	����`an��)�����q<{�_�w](d��a)3��Q�� �!�#눢ڧ���.�cS>;U���v`s��[]���8��O���˓�����c�q0��� �@��_��A�������	2EH��ڤ,zYn�Rf�$������N@����jW��ؤ���jG�A�hhU�?*~�R�0���'�2w�W����[S���a�v��BD���*���������J4V��?�%�O�t������5o<���^mu��EyfQɔ�]�N��$eq�'�gaNR��F7��Oi��N�t��ww�Jߺ�|j*d�8M��^90L����z��1)���~Y��s�W�ւ���kU`�
n-�Bt����VP��N�xRQ�7YT��{EBk�ˑ�ֆ�Y���F�r��*� �2ϳB����)�m�s
@
5���>��4$�oL�̨M����DV
+u��^!� O��d��)�r�r07��B�a�Q�a2yF�uM����+Z�g��f�A�'���j_+Yrx�xo��}L�닏�F4T�&�y�� �]X̚�Z�[�vOlۤ�\���W��n�����*c�E��A�0��T�R��lsr��u�X�"P���q��k)�����s�QD(���� �ɬWW�����Èo-ϯ �AS�e�wa{�Թ������]�Ĥ*�|B]MnQ�{��Y��ى�8�O �+p�L,ʂq�\X:��3�M�,:%_A� ����
�EI���L�*K}3T(à�S����T]_�Q��"2�)���v&FV�X"`Y,�9Q�L�������Nэ��:K�P�<�Q�Y�_c�������DSv�}�]�D�V[��X�{��T��YOQ/�������h`������WT�-�P�J�N�l��9؇Ur�0ޓ��o�9r�n�9_VIJ�A|���V-]��1?@�uZ�>����-�Xm��Vv�x�SO�}3Q��ϕ�g��+M<9� rԎF�;Z���db4�=
�x�2��e ]'v�������h�Fp=����b��(3Ry��?�T'�q滹�Jb���xE����r#��B��s*+��آU��)a�س�V���y;ˋ]0q��"��� .�����+����&T9�W�	�v`Z�o�n����4���M�K8��ţ�L��UJ�����u����8&Wͤ�n��닅��M��i^E�K���oǌ
�t��q���
�K������6�]��a.�vm߄��>Eb�Br�$�^�$��C�
Q�V�S����r���Y
�=!���D�����JBfX.�%`�=[��/���zOʫ��m�տ��-"Y��!&X�"�_6�ڽ)N��y�,�3�Ub��|r�VxO�D���H��g�#z=��Ct���`T�rņ�z���
�&�Ч*�"��c�i���ׯ�����+�a�F������g���C��o�#�a�>��l�@��{m��H�0�j��jhtIvc�A��LNdWJWZ�W���.��\;��BL^�@(�P9,W��CP�2��6��έ/C>�Bk+˕��?I.2��4I��E)��G�i�1%CZ虏��A>��1�r�*���Y������-`|"c R�pY-]�CUts���@�)���l��b
}��E����8�N<w%ϵs�9RGE�}���~F}.z�qV�島b����͵����̷��!�%��2V���X�w#�����Y�	�Ib&"m���ڝg�;1NQ�z�y@��m�w	w��\1��/q����=c+J׉ ��οb�I>��ǻd��7'\�R��~쁞��ݻ�]��^��a*O���E�	l�j���;~��Cz��AV�d�93�68K>!��cQ+k��Jj�|�Smwo�poa獢{��B��e��c��ӷ���*�pL,Z�����l���j����g�h�D� ����G���Ĳ�I�1̂#�z���N����5�����V��2�5�j�a���m*$����!t����W/4�M�i'=�n�*� ��V2��B/��������JWz&^�ڜ��k�6��R?-��f�)��"�D�l���?�EL�^=��I�A���ee~!ږ'�L.C�Hj���a��PT��M��U�l�,mL��'��7��AԸ��#��`�{,�m�Gq�������Ҵ�I�9n"�%�*EM�铭�`z�РUv�s`�-�j(��x���ǽ���T���v���/`1tgx�)Z2o
�|�'P�:��!����M��4s^���uVy=������v��� ��k�-j{����{��$�<Us�"c��Ӓ����VF��VZ!��X�v���D(^�u��+���"��bb�m�����˹m'�fC,=�A���ݓ�EI�n恆1֙�,�@���d���!k� �������ب�G���t:�64�tt�ؐ��=F�o�N��n`[Ұ���J��0Wa|ܸt����^����z�t��JM��W���ұ��?Sԍ�j���uTM�j8��i�'K, ���f�Du����v�E��U����p��B#Ml�L�0M{e�{^F]��^y-f����G�j��rG�:��&(2�*�����_ �%b�vw-VM�Že�G��Q��^���/F�1mH�30��X6}	������ c� �Q���!H��iu�	�j��я:����������IA��{�j���O%�5�kޚ��-M��ڵp�7S��Le�S'��:�;�v:�Nb����`�	��s���N�b�Hp,rG�t��ϒ�I^�z���*��b��oǣ�������m1�u)� �S�>9�6s����Nӏ��5�e^t��b��u!�<V�a��U��~��+�^6C0T�>�Яe������Z}�*��EQ��~�?^ 6h�x�)ZZU )�����h�{���N�!��l<&���wI���l�u��A>~�7l��:D���:%����؄�s���ܲ���9Rʒ��tڶ�fo��*����1�~,��ᴬ��pc��`R��7hrF.VA�/��C�U�N�G���*0F�L��keg]��#��#�gH@a�)Q	
�"^�)�AgP���0.����K��B7E�Z��A�M���w}����p>�s�3�59�rX�H@�]��/#��j�w\�Gf��&�q��B����߼-5��]w̠v)o<��x�`0����%�X�9 �e4��$p��o�K26m5p�)���Qͨ 
&�H�L�#b�ľ���#8|a17.��]K���Dg1pk{��ԁ�0cR�}��fx`k[����#�bO5�s>Ϛ!�#��e���k6��/`�������TQ�bvRE�*s�Iw�%X펆\�xg~�І��/�W1+���W>D�Q��1̞6��D�$o�O �Ϸg���v�@~���#{��%�P<�=1���>�˵��[�u�_i�"1�gw���.��`"�%ņ�
ЗZ9ZA{Y^�Ps�A�!�:�C�<�&T,�c��w��١g���p6�A�m��)��O��% ۥQ魃��砦�xX����fտ��� u�k�W�.M�1Ve,�0�҄�P^���u��ZY>��8}0�����f��_�9��Np��AV�7x�3�;^
F]��&W�+���<���j�̺��Y�dk��L����Ͽ|�PWm�Wt��uz� >�j˂U���Y����1�ӳ�;J��}.�4Ӭ�n�kt�|E�(mdq��*|U,�D���e�)$@U)��r��PY�&񆀕�#�������*���K=,[����O��8[k�%��5�֍Vje��f���䞓���?��/�6���W 霑�u�~[����"u=>����;�Z��?q����u��
Fw��K*�F���]��۟���۸�Yɜ@Lp$���};�C�G�P$6pw	��ّ�0^���Q���W�m�v�"H��N���u�g��"Í!�_0��� `"~���x� ���� �7(vř�mɾzI�؉�h�(�]h?��ll�!��bf�蓠��J�7��@��A9�u[=h�(��B�Tٿ�\UL,t�t��쨳ԣu0�Ż���!�	�
��$�����}�3iB��a�֭�1�v�:b�&ک+YrH|�n�#�F��e/ЩL���Si����3ڴ��?,�l8>W�촢�����m;<"|¡A���<�ս|�UJ�@v���o�(V���9�3\�H2�� v?�G�� 3ٟ���u����e'K��&4I82oFa�$@�$�p�$QOg˒[q�s{�p�;@�r"<�yl��#d�h�+��W�o� 8�� �VUa���o�rit�����z�|������M�Ƌ���.��ⵘ0� 7
8˃�[�o+Wø֠r�+\c�߯-q)��2� �)NG��vH7B��s2�TL���K�L^��0\p�<�N��>�3nd�'&C������1,�aI'�2�)8 y��e�%�F��D�껩?�߭����n��/�ݗ;\JG�^wf_�;��"��,8W.6��>c�Ia*���ښ�,�U�"&>�ɏA��X�k�Y�a�Ź���(V�Q9#ѸI[ʆ�� .G��yeO�s}���k�Z�M������)@B�Mt�uho��v]P����;t'R�n���X~���s:wr�����{:�g\eӭ��O��u�*��'�!j���wȏ۰3q�).��������R�=�
7��j����A��ey����Es���LޱK��L�,/�O19� �}w���%5ίU��Hx���ؕ��
>��~e���+6�r^�v0��'�Wĵ�+c��~FAH5-�t"��V�%i��"�ɨ�TM��Z�fn�T�d�¤S�`ض�{�����%�<N�7��F=���K��}��K��̕�3���R��䁄��m��&eۖm��dJ�����x����p���
ɻBVH���fV�L{qiz��:�{&�Q�8B\-��J�§��f�#N%��qGxi��%_�;�5�nM����t-p�.��b�-�u�8:J�_���j
W �Ȁ��t�����*yC�P�)�Q��?y��Z3a18B�n7TP���Y�S/�	���,�y��X��M���K���ؖz�ڟ��@Ӗu ��'l��E��)��Bܸ�y�(�xk�ț%�
������{0jKXCrS�1��p+��_>:(c,yL��]�CW�f�`1��}�xڧ̳�Zd-Ў���6J��JB��u�4��^خU�"y��@sX&�����z�y��|���ia�f6]�L[���u��8��*d�zN,�hW_R�U܃�P���Q���U�8T���<����RY����B�[&�)XTa�{����n6?�<�'K��"Ć�Ȉ��m� *4�3F�����(>�Y��|�}5d/�W*Q���L���:�A�jN�Ek�	���N�x2P�N9���If�%g�)o�*������> �%I	��q��r���RТ��h�|՝J�>x�@6���p�+&c��e���m��C�霜(2�'����!o�!�.V����v�(Ώ)� d��%/��0" $i����$P�r��뒨�:â��+���h����f�(��.���q��P��Ǘ'����v���N� u�8�Y\r�G��{?kY�F~]�x�}9��a��1��d�eT�{�d��^����Q������i��&�ϧRoN���ei\ ;�c��-�N�AX����(2t2c�7g�g�w"d�r%=n�Z�(<�&���%�˺����ߣU[�(���T. �,3�.�S���������^��>�&Z	~:�_u��e,
'��4���:\K2�7��+��p���!�Ot��6X^�_��T�)��h��Z�KJ�̂�un�;HHa���ob�4�Ĳ&�	fLx۸�(VF��)�~�0�������7	���y�T�C�`��Q�A��Cw�( ��U�v�aH"����3������KP0�\���rA^�ڶ�(-��ص���3�c�G3��?��;xa\�+���Y`��v��
�.�:�i w���Ӱ���j�\��w�Jof�Kqe+׾	��� `o��5K�qR�O�E��E;���HT'�HB�n�dg5�G_� ]�r~��h���Cw�j����y%��W
�hkB�s+p-�>Y1��%~C�C쭝��$�@�\���TCG����8{�K FOyY���g�J�j�#W9�(t9iѻ.g�cV#�no6����y2�#4Z#N+IB@UdK��i�����	Vw"[�P�f�?N	G}�I����$�����-:?�Hܥ��RJ�	]c�Z̧M��bvʊ����Ĭ�	~qI�s����#�6㋏����کR���S���m!�g�WJ纥 �2�Ĕ�4�1�ƫ�=�y������4�L�%��>��)���H.^�r�l���k�}ń�M��6y�Ǖkep��ˁwf^F㶰d�t��5v��M���h(��l\���[�� ^�!��ڦ����M�	�U��q䟘�Q���k�P�%ft]�هM���5�	u������ϫ�Q�@�e���� �������XĜ�!.�:Q���OϤH~@P �>/����e�,u���ۥ�����H�t��HdȢ�x���S(�EޕYd7��,NTV�1A^��T��YT�K_�ڗ�}��؝�h�pm��
�*|E9���T�pr� �Tk$�@���2 @�>��-u�iOcCSU�B^��O��!�!,��I.��ɨ�:����EX*�F�D�VK�02\P�[J,�|]�l��ac\��B�=,�IN�j��p2m�hK����pq�is/���ȯ9#�G�b�7G���Jo2KZ����e�3�4
�[�[w+S0*�V�|R�̝p3���3�w�%���o�zĔ? �ov�c/�����b�C�r�7�U~��'O��_<u�P�������HɈ�qg�>t
fJRnTD�Y�tR��
�@�6X�-�����7h6eJ�Z.��x̪ɋPw�ИT.3�\';��%���qM���o�
;�=��z����A_+�cq��o��P@��
jOˊ���h4�v��V��8m~Q(�6� a�09������U�(d�i0�ˇ����{��0vP�]Q4�XocbşI��<�X�.�NL���#|Bf5_�	����
i). Z�L���:���L��>��(��q�4��!J����v�v�ov�-�e��\4�&M$�X�J�JmӼ{�g��If�����"�3��c���5>a��θF�(8l\���p)|��f��E"5���Ř�����,�^��n����/���FW���5�����g�G�Vx?Xu�mS���\R�!���N�M�����Z�w�/�h!qn�!j�
K�MQ�:H2���=)���<z㶴�*`κ��x�d�o�Mz\�B�ei�����U��7��E0E���ޒ�|�}�cm���l�r��!*��e���� #ˆ�o�����R&4K����43��x��#��t�M�M� �6s����D���K��y�2ʥS�
Z�x�DF���
��jJz�Ӝ?H0#ba�Q�}�7�m��ƪ�й�*cR�V��Vi(i)�����ש|�p�+��Qa@��M�%�`C�xeXMԇ�8��,G�]�2Y������<r�+`�nu#.�\>�A�g�"ą�v�݂^���A�˄�[+p�/ �Ɍj*��a��y���w�Pz�s�܂�H�=&y\�d_A����6�f"{�4dI.�"��q�9��k@�MG�m��c�䕚T�iP����Wh)\^���� \7�gC�xe����������ݗ��̆?�N�ixC�CR�%�XҤL.k�\[�̾	T����������A2T�-Q��)`��^1j��i�a�i�i	j�T�AĘ�%?�=P[���_c�ܾ��qpS�t�D|Q������`V�����%h�&�E�x���:,���g�*N��e�6r������Ms����C�3\��������&r� pPl���7,t�w�OR�eX�(:픚1����&�+$�t3�3ڮBٍƲ�ec�G����N�9�~�(�;�u!`�Ƽ?sJ��W�񼬦�[�Z��Nv���a�K\/!�M�ƽFbC�{~���<c������ 5�Y'�}b��U��1$~�oT���B��2�l=r��b^tY�{Xo<g|]�F��#G~��Y����d�^ʤ�M�����j�/��b���&\��;�����5�c R^��E��SFϹ��ss6T�C�Ewg���v�c�F�U��65���W[�U=�[r�|C	M����y3�v��g�p|d�|�M�Y�N�?�jۿ�-vMo$q�N(�P�g�#�9x�����R�BUw�w@; ��겒4i^� _���쒀c�����hG��2g�kd�2T{���F`�9�窲/\W��In�Z�[�b�njqt��O�<���+��g��f�e1U��vݞ���K����r����G���}��댕�ܺ���R�5oԆ!ҠJyB�6��:��jY9ާ��<�Tޢמ�5�q�"{�+.�/m�X/u?%*Dh|�k? ֲ4���<d�R�t����j�1R�L�E��u���q�{Fo�[�,[�(#}�8W?+,+����;wS��4b����f������7&ߊc����ex�}S�e��.]��|G��i�m]����,�\�@�X�*���v
X��|����=S��p�}l"W�����u a��Pl��n����n��p`���
I�ǚ�۩7��YA��Zj�|�'rr+iEc&ͷX@��g�ɾC�W�����sg�QQu�){�ih���?�QRN��1We��3�̔Z��W�A��S��w�V�-Z�	Q�8�62j��ը��qU����*����>��/F��#�����h�uIqF���E
g��n��(�y�q	l�6B{^�oH��.z���.�X��O�u�L+д�����L�N���?�y��1�K�k��n�owq���G©�_�Z)��7|��]�aA�y�b��y3³�m3[f;_
��Q��ȯ�@�X�J����ra�����o/���hz�w��z�'O���i/l��ӰX�Dc~�J��B�Y��p[�p��ga|*�RsJ����x>��4p81��6��Fi�菩�k,���(�th�r��rbٯ���S���;�^B���\TN�ZO��*� �Fg���D1+d�#ԗ�I�d N���R*յLU�"Ew~��o��>���S4�͒Pn�uD�u[fG�E�e�3�&IM�6�p?�2]e�f%� ���~c��Pʗ�D�`^[��ך�!_` $���ӢGND�h��!��LV�ưw�rS<4��"Ml_4�~gAnv�}�˔Y��,,��V��b������Td~$�f<y����50o-2R5�x.���f�hN��_M0���j�\Y�E����d�O~�p�s��f�^��uFl�z�­,W�ӝ��^�TRWUH�P��7w`+z�QO��lru�j2I�9��L��������Uv*_Ò�L/�Tn)�=<�@�G�&�7��p>�'?
��ݼ_[
4��kΉ�*=A���=����/.("�aF���V�J(6�JK1Kz�B)rץ}&���.��Ct���&��R]��'&X!\�E�=���%�I�E�]�|6�5)��yE�^�������ܰ�sј�\��L�����Z�5+��V)Aa�Ofp��1���ҕ,!���(������:��c�@�+p<K�h�V���j��e�VH/�c�����K$G"�H<T�E�v�P����ڒ�H���!���=���i��4/���L�"Y�V��j����ƹ��K���.nWY����I�~_3�94I�EF�ō�v���T[X�'��S��w�.��Ự�Q�k���idID�RL�U��j��%A�'y]��Hr���/9 ��q ��EEh���	��g�e���������n�抛B�S��濐�S^�oy����@զ_����
gڎ<ܐ�9TӋ�2���ٌ����� �`x������X��	�$�dSP�i:��Ks�6��D##웴7"_�C�&8��l_p;�U!;��m��H��)'�/���e�[S+LΒ�͊�g����o �F�T�Т.=��0w9��1m8f!O��lȭ��V� ��P�)�ڸ3��QRC����Z&�-#�7U���>�Fc4
Mdԯ�/gr�E��_�q�2��~Q���*u��;`�gzQ�o�&�1˖�!1_B����4��ٕ�}t\�q����k��T�!��CO���ң�p�^K����CE}�ϖ�Sq1�.�K�#�Ed ��o�F�nS '��@�d)��<�*����׽I�ʋ�w��(�#���ri�t�<�L�VV�n{ۙ'/��a�o0T�m���MW>�x���?�|~�s:�a�9T��qV�x�e���eԃv�!xP��+W��R�O�R���
��mT�A��[V���<W��D:�g�`?h���¯�-B?5��4p��� �������9%wXU�
�S����9rO'Q�%<��d���;I
������يf>����ffas���}ߐ-��]��
��w")�k��0��řp蛚~�)XKF�g	u-�z�5�U��"5ZFI�d��Q�5�F��2���E�H�mX,R���}������8��c�Q��f�CW��0 �	AB����������I9Z��"�9�;nGs�0,�!"�]Uӏ%�}���*V��YWl�Pt�Y�؊=hiCf����#����ߙ�B�u4稖��f`dwR�ϧ�荄��2��c����s%g�yr��T��N�h���`!���-6ins�T�m��:A佺N���Ub��/-@���>��a�������k��E]��fx�yN�%�~�o�NU�����5�8'ði�鷿��1u����$*��ӣ_$`��XD��H�>ۢ"J-	m�����]ځ4w��՗�<�q@���c������Ԃ�����B��pT9Ռ�nL�,B��A�.��h��3��;+*�ǃ&k���F������
�ӓ���|<�:q1M��X9� a��g�L-��05.f�i���0C������m�p���H�*����|�8G���ɯ���tU����]�a��4ؙ�y�ν| �SA#���`����Ei�Ͽ .����\������I?@L��3�(��N�[{��|��6}}�l#�R��":�mc`eµB߿(Sh<��#sC
�ʉ�/\"���p�P}|V�\�%�C2���vUԑ�=f�Qs�Ր���\�#},c��Z������:X�^�=�
J�8Í�vc���A�O�f�G�%<7;�bޫC窒��z����w"�.��2@��HE9W�J�N����&�#����K��0���h���諡�9P��7*l8XϤ�&�/f͛݃}��&Е~���t�އ�ar�xc�R��.�2��Q���Ћn�?����3⍛V�y�4�(�q[7U��:�}�!펉V#	M�7�e,!na	����#�(��<@)a���:�!���޲?<v!ЉV١$æ&e*�++�3�`xxV�ȑ����V�3)s:y��;�5%<s���W�	А�#�n$�EO�5?A���m��]�d�9y/�-=�/w��]xV�im�?:	'�ȷW}��I2|M�e�`�	�֯kqύ�Մ�Q䠼�M���*���nM<�?J����d���N��\�,��.[��vY>���gr�*���F��#V��u��!;$6 ����/x�BS��8	_Zr�`z��ӭEx�t�Bp�8� :wSAV�7*�%���Zg�4E���*���4�Pܥ��$z�jzº� ��k.���t�Sr�p@h�����6��8��hu�2\؈d�+]v��B�8i��T교A˻��ɂ�Ϝ�+n{��a3;S���՚����u�&��ʳ���9M�� ?`A��Y{�IS}�po�U?�ul�α�;���	��IG<�@��X2��-�9�t�s�l�Y����(�P� ���(���;�1�rTx�7����?���|�/Ԣ)��-�@Ҏ���N���$d[�p@�����:��	_��x�g�w���M�Xn���������/B]Tq+-�B��T76�^�Z����ٴ�f�;���;��X�!���v��2 -�ɇh�Xo�>�:��H����2�L�ׅ(���|ҕ/,u�p�����Y	~��m$��N#�M3�2���u5�4���J4�{���?�u�L��t�����FE׶�.���	�Yw��\��-���B����Uʨi�V��@�l�Ѐ���˯��6�U�����C�<�N���`���S�^�$�?��a$�4#a�c���O� /���W�<������S#�`�-j�qOz����U���O~�¥��Ns�,�e�q5n���it�F5��~�G�>0���н{�T{����ŧC<�7�rɧ�����ɐ0�ּ:K��A��S�� � ���|����Ws�&���X^>n>:�j���υ�S3S��i�F-��)�	���W�����6ʾ"D�\����Y�%��;�Pn=!X��_�Ǣ��n ��V4З�
�i(n�M�-�?�-e�ڴ���#�­&ǩ���m#� �w���٣w�Q�{�=�J�x�Cf��.��)}�]�%�i��v���NӺ��GMe��K���A�?��2��PՁ�	I�"~�>���b���Y��=�-mk ]�~a�y��@��6�����{����"U��ȋ߼(��{]�9���m��0��sRj����Ptc�l\�u��0[�5���w�̇��c�� ެ�"�S�D�e2�d۟���n?��pOֈ�|�>]�b���9��;��d@�k��t��g�D��~���	Ĳ�J�g�.�K5�.#\�5c� ��/ǅ�$�;��r������V��$R~���NK�|IET��l���y��7qŀ�=2��A�9��Ԑ!Jv��Nt`�C�pxf#��zl����	�S5�]}����R�*/���L����N|G��SwX����cU}󭥥��Wpr��V���Y�Yx{����&�v��!��܋:<�y��� D�������5/Cb��?+ʊ?ri����T�Q���>Z�28w�_�����GH-�����␲��b0�D���O1P��,�PXe��{n�|8w�N@SMЬ[ͻ�;yP]�Yn��a��]��դ�7�c�8}�u�CB�+�n�=�#WL=ܕVߗ|jn���C	v�_�,���o�ΐ�E��+5ﱁ������ $e�J��E�pDyFZѣ�������	�P��w�Lp���4~�Ek����"J�6�A5^d�A�����
�&��O_lUL��ڹ&��:>ԃo��^�f�u��\��DS�I[�ot
O��_�'_cQ?C����������&.i\@c�c���)���0��I
5�� ��Ʉ����
�������P�� �`���0��0��g�e�����2_p��*��I�$x݋�aV��k�V#�������mR@��]f'�ϫ��S���鮯#�c��~���	"=˒��ʶ�P��KZ9��ކ�%(!��: E��~.}K� $���0�+&����� �#��S%�!o�� �����9���{W5�Ɛ�n��
-�C��9ј�x�@�_�2�a�+��̯Ί�ioW8q��t1���q
mryM��M���܂�Pj�"���Kh�� �&�����Vg����n�9������CO��<���ĸɈ_���]�&f�	���Lc�%�~��
�SMd�r��f�7�����I�dB��b�	�o>rϟu�1v�ϋ#�ﾘ�8�C�D=y��pq��# w�u����V�?��yࡄ��U�V7�!�dM��Tq%���-V��W��$Ip�%k7@�w�P-��F9�s
	m�_>��';�&��J;0��y�:Q�=� rH�������)$�2\:ީ�[1�-�0�x�.��Ⲝ��<?�f��+��w��Z�@�3��iM<��E��Xv,���ǽ�\��1[�A�K�)c^��fUr�]F}�Ѧ�>����v�qt�>?D��QN��u��r�ߑe�A=T�Ȟ������LI�<�N!f)wi5F!yl��-�<���S��S}%9��p�p��.�uq�Z���Vb�k_"���L�@q���1w�2�%e̍x��C?��?V��\���N� ���|�6��1�h�ǿZ�c�R��������a���z��71�S�Zn����� I�x!��^�"�Y��d��@��J��I"O>0��k���!ӥuMR�b�P��"t��o�*�G� ���-0�lm8S�]�0�j�dEM��|�(���ʷ�I��2�l�t��j���	��2���������ZKEV��(�+��f��f-?�T��$~d�}c��D7U�������Q�|�"�N^�nv�Ǻ}���i{�B�)�;�+�J��f��M)�
0�4��kEQD����@��^����_J���~v�G�K3�T���,��;�4^��˲\0V����Qjk6�v�l	Ƒ0.(-.�N� ��H�3��f�PEaM5c�|�I4�f>w��[�Z`�S�l	�i���h�&K��\�%3٬�����t:;����djqu�(\������Gt�׮�ؚ	���7L6�S�J�@�V��R�{���c9|A��~�r$�j4�o*�N3s<�%`&hDf�fFnQ�ҺCY�Μ�olP# � ^/k�e�2Y���w��V����4�PA�]em��0��\s
�T�k��/�	��V�^�w��.D����$ۥy�E����.M�֋��H�f0������7+�kwo�I��v�?�^���U��B�h�����3c�|���́��Z�����8���
5�s2*Z/}=�^�Ha�!���Y%]�w[='��KS��c���s���Ыx�O�Ӻ��EI�7Aր��fS={�Q#B�E�tv�x�Z��4��	3� �M�o�������/�z��4�KE��t$;�=H¢�Y?�?��io�J:�+9�)�IX��$\�?�)w������).+L����6��v˚N"��v�-�#� �z0Z��ې���F���.��5�d�:�/�H���p��o(2���p�a��~���G������۩�-�Q���
��6�f �;WzΎ�Z/'lWy�������dR�T��|��tyⰓ�����C����𖘯�������ITہ�}�{��_6�z�S�����s�i>��w��k\������n�@��� �Q��a�����L���NY��Y�x����3?�'���k��O���ԅމ�q;Ў��$U�qL����8�	�%��s���s�e0�Z:�+?y�}}Y!UO�K�Ņm�
<3��(���_�0aK���t��3�R����#�Z��"Q6�Q��!4̭��Y.��>|Q�j3��0��c*���ǯ�Hݝ�7|-�i/-B4���9�����ͻ�������h�7V�ʼ,�`V�;{i�z�f�4�T;i�̔eW�����z�"�8�/�����:L�h<["�B.���/1X8�|���jyEx�L⑍=�2p��SӞ����U9�Q`�!�7@���L��ڊ*x��N5Jw �h\��t5�ק�u� ��{6Jp	y���J�Ytb��x�j��1׊Ag`��'��T$c�nR�ĪR�ώK��g��q~�V}���(�?[RV�K��f�����m���>��;��h�
/�={'ԉ�a�ud��IF4;��n�8�}>�� �';R
˟eY�0����}N��9_�~gk)���[6x�S�����jTϢ�Q�718���#.L�G% �l�!�*�c��+���k����!?Y����djxk�5K��^ ��$E
�;UD��7���X(�\dw�;��Q����1ߵ�5���.0S���*�^#ë�� eP�I�?��V������
�<}�y^���aV��jGSӿ���d֏~J�W7y9�Ԡ/�ɟ��G��{����N��e؂k�X�S�m��⪍��/뭔b[e1�;���d�lKL:�x��e[�R;c%O���]���xǚ�1���ٌ?�vb�A'UI*$3ee
�K�BC����^"�Bܱ�n�O8�dw�t)���Q:�^XF�Op1,t�~�y�]Hl�XV4��Q	�����@T,� �v�0V�>'y�2�ZI�m�Z�K1V�e�LV��(=3��upIQ��~�����]��=	%��0 ]˳s��ubv}@�����xj�ږ ��q���!����_�ஒ��p�UB�u�+�O��\z�Sэ�8@ФR#�~�U�F��%ޛ��y�����K�W�D���|ɖM���J���˳�D_(�Y���8��녌�X��5Ǧf��6�0<E��]^Z��ASx�b^��c���#.��!�@a81%$�d��O�ܻ	=����w��i��x>�<�UbeB'@z�D�f����Ijް܃_�}g�F��%��f�[���)ߏ�6@Lz������>����]�ĝ����׏��(�V����`�;�9)P�_!�Ĳ�W�H�Z+�s��g����X�)٩��<F�ĭ�x릐Y��rЂ�m���sxH+_�tl,P��q
����f?�O���P/�[~���뙠ѻn�}��|�!v�`���g6�;��y��2fFH5ZN�ޅ��w,��zp�~s&�3!ڥ�:�|<�͌���]�<�]Ч���p��&���ɖ!r���ƚQ���V����V����Or$�LZ�56�	RYu��=�7�x� ��V���U���a-�q�IPX̻���CsXq��r��0TN:��{�l��H�|ߙ����Eew�.o[����ʡ�l�YЍ�㭐�,�1ޯ-�uBTWpz�V�+�LҰ`����g�Lp��f��p��M��n���p�G���:~\yX �d5ܴ�ІS`߆���v�ȶ�Z����}��^�m�u!M�|G�u�~֣��R1����X�-%����*�5�x� �]A�� ��9,�2��~�������P����EJ]���F�N��ܙ�G�P�m�&�8��yֳ��N�N;�5��A�]�ӑĂ2��"�%z��BcÀ�p���^�ALMe���}O�Ip�*Y�5�yzZ3�����v�"�=���*��Bks���+~ ����T���#Β�x�%-5�G�xq����͂�v\����1ik��^t�[LƆ=Fgl��&��>5~����ظc�g��ք���@BU��{y�<f�b���,��S�$�$� ��3U����z'�g��w�I�}$�o�bh�%�8�Q�+�� y u����|pR�}bo]�~N�ʟEb'��}nDc_�a��,a��u�H�yp�-X���E+�{��]�!3-�6S�Q��E�pd��$!촺�����jh�T`%//5���5��n��ӪUI�b���?�S�����kp|�ь���G��������zw�&~�
:�j��odj5R�r",�-@h�%�u��G)��ʄ$��?*+�'\9fQ
#G1���D�:Dx���P�i��y�kfm��e��3��?n^_��'���#.PAlם/t����,H�z��/�K~)�2{��H����hMZ��$tG'�$
 ����!_c;l���r��Zd���t8E��w�(��8A4����K�� ���u�U����*"�{&�i׍��������%ך��ג��WO���E�C�CD���{�]�j�y��Sê]I�f�n����^=L�1"[C���$�#'Gk�'�!������Ҕy���\~c[�6wǌ��������BR!-mz�p=ѱ�}�������W����\�+�����.&�ހ��Y�|�������bc�q�~I��[��a�v�ڿ!�t�L�r�qj�J�;�N����[8/ҁF�*���_���gN�s�j�S�G:
��T����t�
�>�y7&%i꺺� <������f,�N3���ή�%9�"g�}�L��u�d9t���7�N>�eY���R��������V��@�w�,���d}����<e��0�`mH%��u����M�&I���[KF�V7;X]xKS����^ɘ�i���M"�=��)���L�LB�������J]�*���#����$dJ�H��������q�~���{Z�(�ꠅ*9�t{/�� Et�z���z�i�te]��z�`�ƄH����;F4��?��?�:X�[��j�癃���5��|���%-4�7R�� F�����{�w����B�n��ؐ<N�\�b��
Ѩ��O�^;��R��!���j���L��{$��b�1�gn�t%�m��8��h{����WЎC���_�c��p+����Wa��M�hT7�s@/^H�>�
ː H{�p�w�:
=K�@�H+��rǱq"gPN��>�<�vקЫ]�4����1�s�k�E�#o�Y��B��B�HR�*�ԭr�(�R��O��u'�Qfw���Hs!�K�zO}Uu�hQz$mG�o�qp@4ChO���9¿��AI�}%��:���9��:
^����noɃ� �1m- $����e�	�`ӎ��
q��`_��d��] w�< [�1=ei�9�22��O�|e�%f���e�������8f�� �LHu�,?;@&>�@Z*_�t�ϣ�&}GZ��UC�;N�ů���&cx����XĨQ7�+2�,���K�v��w��4�ͮ�RCą�#�qMX_�K���~�f��H6[V_6�7L��87�a��:��/��Դ7�q���E_ԅ����U���$f��r��V0h�4<"U�?�x)͇[�i���77��_Z�j�����,�D�Dp7K���D�'b�DM1�`�' Rۍ�1y*�77/X�Q!p���EX"Cny�"Ѝ����O
P��WK�N�vS��d0fZ�qg[7�ߖ����9e��Aذ5 ˸�/�rM�ԬG �q&��s�`������݈��8��wpZ��?ݚ��r(��4�m�	k�1�J����	�����9���jW�x��dlj��k���ǧ�<{�@��:ٶw4�>�UUɘ�*�b�((��߭���e��4��[��&�9¿j��yg�;d�K��y���P�=�ӛ	2Ye�U�h���+���o6�����y��'a�v�m�V����'��VPk
�w��v�cE`�M�j-����O���	���4�؉ǆ�L�'��a#�+��4c�|ܘ2��]Ū�aP'E�1�}+<�d�O]�Ӗ���]}G�׸�s5b�r� �Ipo����������۹D�2�Vt����k3Y�����&�^u�˲ރ�{�S#�L�5-�z�~N6�<�&�Y4+��T�4�?*k����x��;G
�4�6<��:P+a�9w���������!7��B���g���o��dQ������ ֔�rB���T��\pp*a}�oż���{�ۚL�'C�ԏ��j{��?m|��GʘS�]����r�Ж4�b¬����u@���F�B���^��7e�8o�+8�[���N��'��0��e��ё���:��.��G�Ҙ/&���E�k�5�³��I[`*��Z�X;ޝ��o�(���£�Ys�gS�A���D�zL��M�gy�(�}��C�؁_a�{,�/1B��5hŘ�ү�'	�@p�~T>R�/�!5#`&��	'C���D�a��/�BG��w?�?�cU��ڰq���`v��N^F��W��]k�@0��v���[��71�P�
:
S�5l�U�΃Ο%�ZL,�(�i|�����oj�ʉ�%nsJgc��$�L߫[v�2�?9���@��Py���y����l�噟�Ni����pY�H~l����*$���4��ux��y�{a!�"�.�K0��t��f�{�������w�Ϥ_�C�	���\k�G2����-�>�B��+r��	����J�K`;D�O�D0Ce7}=���~mY����Cs��D�_��T�C�s9�ˆ�P���R!d:�t�~��1TM^�����(s�骨m��a������m�o}bo�]��n��Ӡ�/��o�	�\�@��l�rU�/���x��1b��`L��t���
/,� �E�7����A�s�aQ�5�ܧܩ8���B���潡�_0��:�j�c]X
�*�9���ϦӷG�/h����5Z�4�Ru-�5>�`����]�1�<��^*&Ca���Dj�YǀV�Fۣ���o�9*�v����(i�a����(�M&��ˎaC�~�ta^��3#�
�&�r�����O�	t�xP���O�5����I~����'�#�Fq������	���tjQ��ze�Jg�.V��qԍX+0j�h.�k����97#����8��e�.�8b%$ݮ�T���L@J�V�l#��ǉ���T�a��el;1Ԥ��-]�M]A���Q�{p�����T0:��Lx����hs�N~|Gir�M.�q�;�0�%�K�Ms�~��L�_�*i�B
����SLָ�W����\�}�D8��z��W�_�OZy8�[�[��O���T
�n%��X���F[l�^
~~R]Hɺ4ܣ�m��	�L�ʮ�z��;�Fr��-(�I�WO�o�kIs�JH�o^�'Wy20:j���B���ߎ؏)���d�Zn����s�+2s�YP�:vcBT&�C$^,���:�C殕�|�6�4��Fc�a=���ⷋ�2��
�穝+��&M'� .��������H�ҿj��3R�xS�����*��Vm�a�ӯfu�W$Ϙ���e�����J�sT�F' M��0
�B��~���V<�?a��i���ܛ���y>�|�H��ER�e�+:L�����6�aXSia���T��x�q�R�1�����߫@~�jv��@�"B����|�O^~�6�8v�/�2��揢hX��
`M����e�ge��o��-��R�r�O�T�WS�@�{���Kv�{�V#���x��*�H�.��EbG0D�ԡ>�r�.�ra�s=~O����ߏ�4��Xd^ǭ:Q��n� v���Nw�3�X��`��"�(7Hi��#���+��-
���y9�~H��$6$�N�ɞE��y�W�~^�����_���f��&�p�AP�mt\s��9��(�I=�����2�hWyKۋH�hGގi�,�=�?T���{)��VQn��D�AϬ��vp�2}�+���6HUV����uoXv�9�
��Ki�\B�\���	�����G�q��ֆ
6P��Ʉ�a,G7���l-$�oV?��?=�f�W������b�r5�q|+`h�8=��|r�#�}j�A�;�p�]=&J&�d�����_���M<VD���%��hp$�Emg�F�R��}b�&ɶ��X���bb,l�=l�)8�L��ʢ8�w��}��O9�P?���u鴤>0h��|i��<�`c�>-J}��v"S~���@��[�2Pj��A���2_�U:3TA
���~k�����4�K�ΏvH�Q�e"�m��N.'��مC���2�����9{��p�Z�C\ƒ�zZۻϵ�Ci��!�i8�Z�Iz��'ֽ�����'
ξ���u�+H&&�{!��X�kwC�E�a�L*��0�ѭ�g�1�+��t9<�{@kU	�Pd��.��}x�-�E���|�e�H6yo�'(H\a��\�p<;��CR�SJ'��*L���X��Fi��s�����N�k�淨��C)��f�2�9��Ӵ]F�:���^~i��~��%w��O����DWw�#︤��fEI���#[Ȋ��x��tF����t�jz����Nډܺ+Ypi����(/K�(a�#�7���3tR*��{v��M��u�M5/��6����X�h���Y����`�>HM�Ԍ}����-�I��ah�c,Cy����ى��5�ܻ��L(����JSg�Y3�/�Mp0 |�f\�D7{����(���rl�u�t�6t�) #������`�����OU�d}}�S!K��O�{��n1rf9����Nu�p: �J�rŷ_W�w7�{��9�'��{�Q�� Ś��&�A�O]r�t�-����V%Ψ��d�4��~���)>С�E O]γZ�@]:
t7�VZj�0�4^����Io�
?����=8wR��z�كs_y<��}�7$�OC��+'�.�%8'���T��p�.�8�I�89�м�K�<������?�7
��&��#\�Q�GWL
�u:�VV0�*�.��&ѕ�'9�򋉜T�*�0b�kU��xa.��Il��b���؍S���U�pbK�,ͧp���t͵�A�t�JD�i�:�pAz�����8.����`>}�ς#�C�{���D�M�r�n�Rb{��%'|�as�y�2��,����1�Rk+s}B�Y�=ȯ���٨C���Ε*���-�0Q�;�6��C�d�\hx���3��i'�И�g��B�bM�P�6^��hy��:������>`�9`T�""��e��k�!��rl�s;؅���``y42��!|e.��`�?`��J�ʟ��ܗ�$%>�1�'.��Yb��#�����]�yV��_,��vG���0��ѻt;��󟛲C���F@[iX��å������7v�Y`����wq��:�6�3��|�$~����V%���#
���Å��%�2��*�v?L��
S�O�˽˺��s���}q����\��s绱$��X-�X�n�&������O�=8���πt�- �b��;j�G��_�Yh��3��ol`)�S�mH}q/�ԑ��+��4s�?�ɋ�#z�	|��
�����v�w�ٔt���U��߱sd7��h�Λk9
~�D��㢕~vf�MD���X{��9Wd������6c���B�<,�R_f�K�)���������'_)NŨ4s���ƮN�m�Z���E�*xܦ���Vz�S{9��]�����l��j���[EFĲw
�y�~�P��$GZ����_�����K��^A�]Ѭ�#3J���4�ʛ�(Q,[�s��@uf���\&>'1S�]|�Ny]+����s���������q�kT�M�RU�Z|#��6�i��bń����J#Ca�ܙ-逇<���rj�T��q�&t59����'�4�e�i9��?�y���V�.;���7,.%�� &�L�5��x��O&ѕu�O�x���.� �.w8��dǣZwP�1XNO������U��ٓ���I%|���:|�=�8�Qp�
��R±�x{8@(��bE����~5v���c�/��c��	�ƅ"Ӑ�����m�d$�>��  |���B�Ss�7NZ���N�1(���N��\���Z˘v�k�T�`�6��s�*��3�P=9�Ld�C���p^��i�:x���zb{�$Q��یê�̷\��Bܽ�c��R������_���*w�e&S�����\��d]~�ps�]|��rm!9�H��IzL�ަ�,�I�^�4���L�݄�7I�W
F�-6�4`{T�V0`�/Y��+��-�p<ɤ:\{��md���[�n��W�E�!&FAh1��bəq�'�&�&`)�Jh��U���^^&^�0�P�zR-��x���ݑ�.��`�H>���|o��~�Wg�"oj[����vw����������%��,k�I�B���8�@u��!��J��I�xf�������n;~�~h�N/�Xh*����3z�Ge�����+���������g[��ss1
"·t"A5�+iϚ�'X��^��+�&x���E�"�4�t:L}� лwתd�nq�jlc�����-�D�K�b���'��XG���g�5�:s%;�?�k��9G�aw��E�}��KH�X5�C�$��(�"�u/{�wh 3�j֓o� �430�Li�ǔ�����<��d���cR���X�?A7b�^�#�5u�͸)� Lo�����p�k�~��S�0�>��6�Fy��֓� � 7��6�w��ޝ����Y �<N��������̧=�"��@�_��^1���?�|�P�	�1�x%>hp��~�03���hy�%ŀ�^ED�[>�dհA��x��;cd��yH�������j���eq@�C�߈�������F�!@}�u�3#��GCdy<�Qv�p�T)���*?ս@`� ���K �ݼ&z��	'WR�J�{5�isH\��k2Bq�E�O�ƍxE�w�ݻb����8�a�$���D�n��j��('4��>�]�ϗ߼���w�?�ET�j����1Wì@wߊ�;8L�L��_��}d��ab0�#wTm��n���G5NF��l
<��0����d�Ȭ�q��	n��	��+mF��u�_�ˑ��X��5�&4�}�������v��Ț�5^��Pa�MK��^)!D�y��Ƈ��=]�""�u�\(p�n�"t���{�v�\ ���S��g*��q����U��B�����%ȟ怭���_o���v�6��Q�o�*�L8��Q�V�+�S|�s�$ދ���	��|�䌬#]�3��7CW#^K��87H����"$��_�\��;��@�jX=��g
u�L	���$�pKQ|x�*�[�zL�� ���b,	۬j��o�B;����@��3U@3��}m�XDd��3�3ݲ*aF""3^U�7b݄����~�{�v��W�kӢ"]C�!J�W��񈔧��e����X4�y.F�#�o�#�+L%��4M2N�1�UEE9�n��㭃�{!ň;�`4���x�,ֳ�%�>޲?��F����^ɗ�0�m�l�_�}�n&N�*rO�h�H"�ĺ�ʎj�Rm����ᚄ��u�U|�1�-��8��-6���Τ�5�[!k�O"
Fm�/��m�~���vc �%e=-�%��QRX��:]햎x�pw^�̩�� <�T8R��=�^w�Q��:����彸M�K �hl�@M��gK�g@p��Tu,��N��I4k�m@�kE%ڻѹN��=�������x���e�Q���.h��Ao��К�in`�1�{� +��K��Ѝ�p��z/�g�Z�=������a���`tA3|(�?���wrO�L�u�J��h�����(Ս�~W��_�@��{���#�n]�� i��`��Q���jU�z�U�͋ȭъ��Ŋ�������ʎ�^�R��?�,%w#YH-ߩ���]O��S���ta[�WQh����tz�u� չ
N�8�n�eo���C�S	A��ğׄ�>��D��s��c��b�}���T��Z,JI��iT����.�_s'�%�/�2eЗB=�q��i'��N&"",k�:��̩\\|[,�9B����.5l[g�� ��a�yF��g��{Ũ,3�9^�Q`.Q�Ŷ°	),����7O�I>�^M�8� ��j�-� �rp���W�\�7qzW��7��d(���	O��i�(�rH����xFe�Ϋ08}!�v�N�;�l�6)�ia�T,qI�k��K��O�&@��&����Qx0��u�͠� |:�~g����r�-��MHk-_������P�����v�h���숗���-h$�_`�6N=p<t���ζ-�򽛍Oxx<���I)�2��5�5�]��_M��|�p�r�!���ʒ�^J�լv�*��cm��l�<��S��M�4|o���_EV�f�OA�]X�XE�ZO���(Y�q�M��+��rQFua�#�է�1�60dor�撞+BS�r�D5'A�5�L����7��M��?����|������9l���j(�?�P�F���x&܊��1�ef �����Ɍy���	%����ˍ5c���+�^�C}4�bŦgD��s�l�q��c�_(�=���P_�_y�$*���ڨ1U$8*s�� V�'MLo�t����W���2���!޶t�˶��bz�����#{Կ��W��߂�h/o �r_^�/w����O|���g�ĒJG>Y2reF�Z�C.�t�
�/�)5N����b sùF��y]�R��.�X3�d��g�����h�����*ӧ�>xc*3��R�/wf���v�����������1�����ً �٪��k�5����t?�Y򖐚�F�j�_#�)"R��΂퍽gK�����A�zv��Iq�|���z&��i�	���B�h^��8�N��tQ���\����,��>��7 \��F�|)����WoOr���7��=���4�!=����Iz7��&'��&EB�۟��Z�Ȯ��i�*�A6�L���l]�(�����B
A�)o���aO�/=���#K*�Z��<��+쓮°�K���a�� ��?m��*�����`��vM G�xq���vG��H��C��	
֠c����K@SF���'���ڗ��Mn'R{�O2�g��;Ox��|>�Iu�o�G�t�K���ed�A���UQ�M�Z�@��75]�(�����s��*1'��ЂZ�+�$0a��2�D%���Ǘ��C��u��R{k�����,X��E��ᬽsVb�*QIiq*ɐK�p�hL��7@�`��Iۦj���3~�`���ͪ���/��Dox�12*R<��T�Oȗ��m��-*���z��m �)�/j��uG������v� ��Skf�g��*��W*�#F�EV���<>Ҷ��Q���A|xLIk�w�r�����
��}k���{G�=�9�"��P=<�<�t!^F3���qHa���!�AC��PY�A���<W�����-�af�O��Z�%I߂G��k�H��"�oӕX�:ή!]u��fx@�E��q��N^Ob`�n��w��e��!	J�j�HVH�@e�9�f<�3��y5j����.�ů�+x�/F�����	� S3o�qnޅ[�3�a�E�"3]�Q0F:�N��Y����!'/͎�����p����b?>~a�ibh�@�ؤG2�H�T�l}mH�N�ŏ���F�g�Eh��`c�zVɀ���=�x����������٫�~O1�e0��l��y>�j\F�#�H�vb=�1q�q�6���_t<��7�I��[���.�=l���L�@Z�#X]�3�՛2���r�j�}[)1M�֌�
�S��=� ��С���Cx��Q�8V��(%4O������͹�@�oO� �&��eg��Lmgj+���P�VY�kh�XL]��y "����2C٭������������0��tuP�*�A�R�F:z�C�#wT�>�g��W6<�	�!k�	=>�e��/�W�����#%Z�g�%��[Q�zבw<s���.ʸ��5�j�y�>����Od�I���2���hk7[��������j1�g�e~�0�}`U�����{��Z�X�Y\L���Ծ�$�>����Ԓ��;������h��yS�=c(ٺZ /3��k �q1}���Z���NJ5�H'`B7�'nG�f޸�� T�(|~5@ZGx��mG֎��^���Jvw#@E������z��#S4�_�K
��ԅ�O.�9�0*���Z~T=�b4c�1r�^�F���"�crT�Ns�N:��^F�=�6@"n�ϴ�������հ�����h�H*�\�qᅙ!�S�
2�}����	����%^~��D�8�=z�N�T�I6>zP�_�fi%*��ܑ�<��
��OBZ��p��,A��>��H 
��x�Fq,luO3ya<��g94n���D�8���=#�����b���KU�������\b;�]��L�H�#D�ļ��+6��as��X��t�;�F�)�(A���H�����%,x�'�`ݴ�����Y�F6H7��>�^�i���XL���.�������� ǣ�.�Q�#���� &L�{Ȅ	��b80;XEEf�AO�4~X:mcH?[xe[����A�5c�{�.���Ģ�	��gr2�ae�'�
�f�HE��7��1�[�@�KU�q����a�} ��9s��m���T�^��$�"���V���� ��$�}���=��_]٫�~}4;�]��-��90�,������UYw�����q&ܹ�2|J���=F|ި�b-�$!4'>�����g��ҩǟF���~�i��B���xp�9�Ch�qEQ�+�NvU�OI8,P6f)\?I�}ۋ-!���d�� ~PJ���2e� ���_�/Y�/���X��g?W���k�a|<�,O��?�<\��v�N�dbVj|Ey�EH�����U[������Q��!�B�}L9�#��sU:�k��I���We��G{��k�N6�y��I׻(�r�F@��n9�:�˗���1��7gb�W�F7����_^�Ӟ��({t;w�U�s�t�#��I�=L
����O��L�T�jBZ-���FV,fL�U��g��|$%ar����[�:�՗�W��[�Μ�P�
׌u$�$���Y�{~4��dD0�ؿY6����0v���U�����_� �8ט����^���eq6����u����:\��=&ێ�#O� ן���%� ��ML�S|���}t�:���Y�.|*�+�bgA3_���G����:w�;Z�6�>U.����wۨ����B�D���H��c�J}�sT
�����-���Z���N� X,0�w��^AȻ�/|�_Z�O��7���ZT� ��^��B��+��?x�54���r��3�. ��<t���W����bg� 0�޳l$w&
oz�2�
�o��1��G�h����2bw�&��Hh�x�A��Z)���$د�u���{$��[�D4�~a����4|ʯnfNz,3�8,��Npm�^N�9ٖ�Ї-�?,Bp�0�C�
_��/����9m�3su��.���k�\%�7x�
�K���k���|P
����R�?E{~�ހ))�wO�?�/{�B��DD��2.7
C�愃��߻��;�U�{�d�<� oaAY����T��x����D�f��Z�C�7��8��̠��7�r��}&X���d���6\o,A%j��Y�U�c;�r��n~V0)��d�-�x1)�l�\�dq��+&MQ��J�i����x��n˱���O���k����/>�������,�� �ba6���j��pYl�hM�-���L� G��]�vH��+�~''^U��Fe��kq2	k���*q�!��n;�Z���$�aR�]��~\є�8	����B �2���u�z~�q���q}�x� "v���_��v��^�����Q,6� �nW'S��/`�$���B�_�<y��m�d4����]{�X�X�-����L8 ��mg_��ޏ	X��a�"��P�ѕ=�%@��%G��i���+���cMR"-�9��D���&��������1h� '�\m[O�:d�G��d�+�ࡸ�mY�9��3|�*�⨑OR��T$�$7L:P�"���2��j����� �a>^���Y����&\��������s��o���7-	�u�c�R�?����7�z|�pYm�g�b	�E�RB�co�Ka��F�*B�i�t/��t�����"K-9�F�@�_�D�!ӏ���,��Y�/ۈHP�ț){vf���1-�>���pht�r�&�
�4�rh��&?� �H�\�>�{��p%���)��/bD.눬;}�G�,�4��(lX:�Bu!6:}�L�tj�y~�
h��d��-�3��9!�Ư�^U�Z��G�ƭ&6N�a��vK�d��(���M���@Qߨ7�� ���q2{ʔ�)�k7�͹�yp �ڰ��������3��1YO'��XH4�?�v?]GFN
��>W��z�Be���+t�"z�L�����b����X
��FC�V-��yn?&�e�v�Bv�g=2�����]vFt7�Qw����<���X���y�? ���|.�!l-�ap*��5�{��uyv�d�@٬�g_0����/�!��LT��U�tlol )ן_�o��sΌ�5�t��92>����~:!�t��µƮ�D���0�x����A
�ָ��0ӹ˿}9�_A�Йj�����^��:t�;���O��H���eDtJ��ոx^z
��~(�w����g��E��ڻW����g��Lgj�UU�?|@ԝ�t4����ISU���p^�uxY�qm�~ܸg��n����Wjt����z�� ��	$T�%��Z-��?�O΍D^]psW��qgNE9�"�b���la�Ũ��F����e�l�0�fAe�;p*�=�^�Scj�#�qި��oFlg��+d�] :s�o԰y1 ��r��z:'=G�`��a����)=�� o�l{c�J�_Ɔ����~~E]�u���t�Z�X�|)w�dGJ����F�z�1٦~�cF(��#�;ћ�{B�Hk��0#B}��٭�;	�q�8�x���Z�Tc���3��-�|(d�].-h�W]�y�1���b�\�4�Pq�Z��*S�Jӆ�r	c��?��$܊�G�ؓ!��xFm�_�g̾�cP1����*6Q�$��-r�Z,2�	4- ��U��`�*�@��D|��������zc��>�еS�-�Z��	?[��	$�-��.�Y�SHy��wB�x +���wvGS9�����\m.��Hµ���2�1�}s<���#���&'/�����g��F���`���[e��}wqB"�΋�,��k�JD���t���CѨ��׼��J��A �܆�(6$��+���AfJˎ��|=J`*������	6*^Ċ��^5[�Gg�_�̌u��I�=Ɇ�P�>���o�C;#����2����Ԇy���ʆ�$������
�/�=3�9:$�p�~&+}2A`Nc���`���?�+9.����@�:��ޢ��A���� ��*Bno ��P�r����s�$�g�5l˯h{�1p��7&��E����[���b�1�y�.a������@}�&	��/c�\���T�ۢ�|Ölg]��l�+�/��M�ho�R�mKă�7��3�G*�{zJ/������1vo�L�Y�[�j�{�?TDDj��-���	�,�n��o��u&���(D�<v������o��]궄�,��8�[O��E�-�E����0-�[t�O�_���]u�#*����M
�p�%:�:�їԞ� ��j�G;��K�!w-��C�䜷Ϗ?Y:N $��8M��N����r.M�soGM�kj�^�N��Z�x�UN̛hk�@���&�P"�Y�Rߢ�wִ�&پ���\7�������)H�v譴���	q�什�E,�s���j��{�ĥJ�z*��{��D:6�������}�����]oR\���oԝ���g�i������OBd=�Z�q�uI�\ఠui�����OK/�j��R��u4)	�'G�`��yP�(�����ň½��5W[�s�L�+�b�$lėg_��� \����x��wFR�����\����ǝ�|�>�Tc�n6s5��]A�B�p��^�m�J'���Uf��v�X���Ѻ}��d ��`���;F)?=�ԋ�ʟ��i/��A韬��L4|Q�,�l�_QD���s�h�_,��5�b��]�y��y�1[�RǶ��}DZ�d�9�ޣ]���S+ʃ6�ܴ3�&��9�,�d��H ;@�-M�E�A˚b�1�
M�D>���Teʛ��Ym��[���i\@Ir��]8�j|���:��;P����`~���#�ٯc����J��T9k��p]������7>ף��1(�h����!�Ղ#7�}�¬�^y�n�Zw7�����K����B�K�7,���HCx_��5I���kT-6T���n�#�.�gOZ�����Mw���ܙF���`�!�h԰�b�f����F�H=k�]���c��W5�q�y��g{`���e7���6	�`bՋ֯e�Z���m�����2>��Hj�=�u��Тs���]9HA'��۴��ZN�j��� `�l�A�u�4�	Q
,�������&��V�?1�8A������\ڋ%W��/Bi��W�C2��t\��2�+x�,R��V�dp8+����H�>�Y��j$LncƏ�iٗ�CP�ɵe#���`���'&0%I6�A�FD���nF	�`��v2���l��<Ӣ��'�ZR�1��߃i�~�ݼE�P���e��[�� C )��1�/؀f��b�>�mY���S�seiQ\H5E\�Z�$}��J2\!�͟;�I��k����NF:o|�A�f�Di���@5��l�.���"
ş�ed��	����d� c&�F����4Gyf�j"�j��PU�:A�����h����R���{J�0l�VĮw�Х�iēqCr��}G\_��/�5v(�������1JS:1�l�kg��yQ[���r3�缮��`3�f�]<�{�j�J,�O�Be���e)Vh�k��?r
?���]}��|�<)[�5�q)z�[�������Kl��<�5u��8Y�Z�_tc�Zv}��~�}Gk�fp�K*՞��������"V�)>�)�q�i��R�n'��fU��Q;O,����<�v��w�O|���q\7���4fyK����ϩNUV������.�聪c����} KQ�1���n��a������8�{�S�?��}2�� i�5
;u;�f��g6�q�����Z�&��x�bt`PO�Z�,���X�݅�~W���N<Y�5����)(�~�����=���4}�-q�X���MpUV�P��,\��._E݁)+��������j�,�g�D���2��T].f�G��}�p泭k���wR�>� �ѨeܢD׆7[������OwT������&H�_�Wi���� ����=v;7vq�B����w �@y�a(�4�Z�?Fga�����^�y��^�M�K��ٱ�kW6�����g�.S j_4=��ĝ���Z��Չ�B�IfC��x����Jn��\Y�y`�d:E˴ �ԋ�n��1�����qr�	L�u'2*ɿ٦��ِL;GH��(���0��J��C�"�W&P�;�R.%{��>�g��%��'�B�	)�~U����k�h�C�X�ӑ]c`X~&�q���r��;�k��i8Z������?��͞C� �yaA��5�ӷ$�k"���8�r�����dV��8��T~���ZXA���yA^�,�#"�(7�Y�ueo_e�sYT�S#Ty�6E?jӣ���E?��G�ix>4\��{酎6%U��&Og�(z4�P��7��1m�d�Ue��	h9�/
^�E��:�%������pje'M;��ࣳ��}؈��!`�a��_�FWZ�B ��IER�E���|�d¨.�7�7��X�F�ٺ�|y�bѲm����0]Rdۚ�B�: ��{�;�V.��w�m�٬EE0�л�t�x�:z�\�h��QM��(��&5�;�m��F��xP婌^Ό��؋����2\�,旤-�d��$�o1����jH�����栣�ݞ�{��BN�b��s�։�ԓ��� ��L]�˴�hVʎo��5��3����������.�ub�=�[(�m���q��P̹#�Ogf�����уt�d1���汈���YT��5׳]�;�*Zc��b��H����)Ԯ�/�.���l�� 7AA��}U$u�}���H��o�5�K�m-�,�)�0N,��������7�]<`o$���p���Q.�=]\H�%븣7|>�Q��Ǉs��=�u���A~u:�/�m��C�d��Iځ�*�fro����iQǶ��m����i�NS�74G�"eZ��-�4�Ԥ4���_k��9�G��'{�#w�x3��"�ݲ�"bm���I۰q��]Y��K�G��_��H��Ue��Q���� /־��݅�y�������C\>&��W����I����c\��P�lo�8P�zl�As)a�"��r�+%V#�����0��{B���tZ��7� ��_VM�B�DeB �yrX��E�-2_Q�G����d����P��I�*�f,�����`PRȿ�O�����8��)�	�C�qV�"Hτ=�� ��0���˦�R?5�cR�:_�i��p)��v*�����RM"r!o=oO˳�k��}�d���W��#O��-���� I��Q��I��L{�Kt �b7&�Z�x.���wK�m? �@jP���C/�v�B��L���h�CĐ�����CQͦ�K�\���J�'R,h�L��X��+������3��S�Y�q�D������+�d�eTܥg�4��2_�T\e�?���e��1w爦��<ϲ"�6�_�,�Q���>s��m�� -�S����k��uK����t��Xl�ߤ��9{�\#AO	v
vbD���(��fu���7��ڳ_9�Z�M���(;��<kl�c�=O�M��4t�����GUsf0n��7�H���|k�"T��cY�BV��u"t���f��	>?X��kX���vRf����5ua�"�/�6�驐s>��� �Ř���{������d<�=x<�ǚ�Uzo��][�%�%�ێp1��'�m�p؆aJF^�|�οs�TQ�2R�?����C�=!��6-,7�O���,sZ��=c��UG�P��L�]�2�v<0x�;*�tTr"���	�����ѩ��&=)���'ڍG1n��cfL� ��^���HI�Ū�K���B5�_�l �;��:���b�����2�<�[FX����:<�A��� �> ��p^Ijڊ��=ݵܮ�+���/Ԁ�zf6�wU٨G�d|�Oi�d�ؖShxBjBh��^���X1�Bj�lcl��JEl��Q�|_�]�����eT��;�}��"B���-}U�_�L ��Q�8��w�w*�n]��m.U�2��ۯ�U	�MP�*ǽ�9��vU�f�'���)k�äĐWŴ� �ź1{6�I����u�{Z��,���F������]�x������D=aM"�^mWh��N��;)<zσʀs(n�z�1߇��ٖ7`j���ڛ�9����#"ܴ��̄���q1���P�V�X��������P8�#��Jqw��\����81��Y��]
�Yи��|��E�[�G�y-8��pO��F�km��(Lk��N,c�Ο٠%=��4,�,yw�`	$7�-��oa��{"D�D�����\}tG����,�a��2����ޒ����3r�ƅ>CP0����LF���=*ʏ
{/��|iT�w|�`��H�����׷���`U��:x�G�&�쪸�u��I�ؖ������B�ޑ�G��A;_)Q%mm������
g<d2���)�N���o���r'˹�6y�8�B̓S]�ǡM��n���Mq��}SR�4Y�E>$g�R�*�%�^�G��/ωn�,����$*���uQ�	�gM�ps�j�i��jǪɾۤ�PP��-�v�@�H+���YS	�l�u秇����G�L����;�e���{���'�.�.��(c���8z�2�6�
�Q�����^xlR�۔u�`)�Z��p�yvx����4��)z'r�1OĚ;�#�=	��b�kra��Ӹ���u �el��ˈ	_&i�~��`��#���zr6�����K�#�ɛ�ȝӒ+�[�"M{]*ޡ�;M�.��!ο�Ƅ|�f��E�鶭��m��`z��jC�*���+�_���Q�(҄����%�:ӻL�pQ�:��V抖�6J��wW.*-�J�%J3޽	3�OqP�-�sFh+�[��F��O��LGh�����N��
g���7�D�)�Й�� �+�R���bg\(k�M���ss��*m&�jC�����%҆�y�����7��Ƕ5\%0�r���PV�)���C���f��v�Z|��� ]0WR�@��%�N3�I5[0��ES%xo�P�Ý�[*Y%��XlF�/�㼔�s�b$�^P=���л?� <N�;'=�&}s���0�0>��7����ա얉�]o��_�a���� |^�kl1 �pw|�ho����������v�:��`������hu�^||�<1���g�
dO��צ$(�h%cY
R�8HJ�5��Tm�L�̯?��v 1ݦ�sC�;l\&�6!���,q�7Ց~��c}-�Z���f �@�����Y�:c�>>�Ft����=�m�ɾqMg.P��@a�pz� [�BM�����r���c�Cd�/�E���h���1�# ��v�up?"�Ǡs�`��&��͂�8Ѱ���*���$�eR���㶟��f�,���7(��ˤ���$�z���:��/�ԷҺt>��`B��Vjde���A�V��o�zA�'���'ߩ��g��ZC=��ѱ���0Σ|��8��A��\�e����m�}�@��3Z�^��M�t9X~�Oǳ�(`�k���y��RL�~&��M�p̻�h�40�f����a��'�[�;��Z��˂:�b��Ѕl�:�$�&���k����CԂ3���I��
)!bY>�}կ�>����n5��UR ��T���#/q��p�y��4����*X��H���/�+�0c��|]bHm���}�mӀ毟��"�>Y�jW'V�t�� �8*Bޏ�{�<�C�E'�:� �!��F-ן����t5;����
HI_��Ĝ#|�#r\�ق�}:��������b���T�}����#&3��
����c��/r_�	a޴ի��R��l�^�|Ĥ����DF��n�	��^��e�m�����b�Z�dq���W�G1�RqqLB�`�"a�6����U�:T��.m+oNf�:�>���z�������CU�L���/#���X�R���X���e[](��N�RY�{(���چ���[�Aͳ��3�4P�����<���H(��cZ�f@i�����q͔�,��]�Є{�?X�m��bo&k�@T��[���f��N�/mڏ<θ�k/6#��m�f �$p��KIl��ĝJ�R�0�����,�h��@�W�SqrJz��cA�UC]��t��T|��w�M�y�=�_��7�����%?�.�[w�����\k�T�ra���ˤa6��h�7�E�㕩15F�?mg^��ϒ�#�C�e�K;�I��h��0�N\��L�͌h:�/(g�G�r���"*8<�MY��G�)�q����s��BvTxF��V��P�<�pgEZ�E�t~x!��;�R����d�6ߠY�n?'��x��lr�Ljk�{b��
GW�wS'4��b�kTy��GB����_�ႆV#R���m����B""6�U��S82�-SkyAO[.�)��ם14��?��e���d�Fc���㻛[k�*E�P���.����-}m�^Ω���N�r�¨�{�n�ǉ�^;�����u�@�K�D�AT�q��i���R���gB��r����UD
5"���MC����Es������'iO��V�|��e3���#�W[Gh�mb,	�[��&��Ki:���I�/L��H��V���́����L� v>ե�G�����ZD�%�^�;(N���3��`$i�������UC��l�d��ф�:�y�'�@'E��:�����������z�p#�*��\ܥϜ(3�����Z
(<o1��Es�0��I$��](l����������g�� P�v	 �k�p�PL��J����҅mn�e��ے��Ҍx��0��o'zʐr���-��Ew�2�}�PϤ�.�t�F��q7���աK��)���-V�p�]E��۴��L��2k�5��B�E�#�T�乍>��yT��9L���	O�zf���U�+<fw�i���O�y��'ZX	�r�P�A��GpB�}s���Cȝ��JX��	�<��}1��S�?���½�Fԁ����7;�r$���<�u�B��0�Ǚ֦�t�e/$^�� ��zȹ~�[:�3?sU͕$��v�n:�|if���=��a���6rF�_V����܅Ǽ5��l���|��r�v���ǬvW��v�$[S
2�nfː�k����I�Q��RRm�2�|T#nպ�E#��)�'K Ь������Ժ<r^�c�Pwv7pg
���[�����+�r��QNȸ����c�;�0��tO�F�Q���}˹1Rsai�O�榀P�M�4���O��'{��Yw�s�rƴd�Ý��P��_ai�0q�o;,�8'��u.x�0�#�ЪB��F<Tv��}�-�i`�^Q��K@�`�5��vmº�P��5khsD�79ZƵgQodz�ȫ��s�AC�������J��F������2bq��k�#���� F�W��^vp��B��*��+s� ��y�d�M�����1"�8�?��xͳm�uށ�<�Y��0����̽;�����1}4N���2wq4h�w$�8�BW*k1��yR�����g�4AS�cV8�q�}�eXpp�%/0V���G����z3�t��!	U'W�޲�F�$�J�_��5�׎O��w���φ����%ҷ|���VR�%OK6�>[˘�R�o�Ugt�Xm���`���4��4�E��m	�'x���)ۦ����ßX������
� �����Տ�w��_r�z"<Q�+��f̕�Y���-L	�������:��ERmG�����A(�E����o�]�C8��C��d�3�cr�%�v��Hey�@rC�t�RǙTa�^Y+���PR���=�o��}Ց��R���n(�Ե��x�؅jAe�G �!��P�3�� L�
/	}B��t\�R��I=��V�q�sKi�̩������D`8
��%�#�{n#6��X�T�
�����b�������^��`k�LQq�E@%�וVگ���/�0�PT��bf-}���5k5z�����.Yl�	��{>�ɬ�2��*W�,
�CB�)a՛1�ԚoX:���<
��Ks�m����U��9btA.��e��� wb��ñ�˒�$�B Z5���� ����{�Y!\��B�*bFKʧn(�[=	�DM�+�'s�.>��G�����@.f�!��\�,�������5|���DƑ>�1<v+rN�����Zk�ʲ7O��{2 v��FA\8/rI�T���*zq�NS�+��yi���wq��XEvS�4�2�D��K#t(1?/J�5j���O`7�����R͟ k��6X��)����/%H0�LsauP�ܑ4�4C��97ڠP���c�� 8*'K�W�� ����C��d5>���,�#���M:Z��P@c��|��v�k�;��渟��B-g�pw���3\����bWX���$��5u]~	d����]3�(15��ȁ�
�A(`w;�DS���l��:3��E���CP�boǼ�۬�	!rT���)�%q���H��l�/H�A�6mU�,�����B��<x�c`��D(q��8���4#1�rc��f�� n�5�C����+���z��_-����ք{�����w#V�F|���p����.Q���
T�7c����fq3I�#��D�f�bA�C�P	�F�4�I;�/]6�f�'���N�@_m2�؇m"��W>/J���N��Y/`Ԭ!�"�Lm��i����Eg�r��"�:r��i
ÓK�m�f��RqՉr��"_�/GY7�rq9p��`o4��% -.4�Ш���B�'�):Z!�E���0�c?����)��@�90K�ӓ��$x�I���˿p�ݸ�HE�N]�m�Fe*'+Rp�a��*�F��Q1U�F7��J:kHiHO��h�P����boٻ��n�a�,�eoa[}?�F��GZ=0^�Þ`���P9h���8ڐ1=eƾWـ��iE~�
��*6�fj��!�3Q����2�3ņd��2��iLT�@Ƀ������aV솥�ޑ,G�[���CBG�訤-f{���8�A��1�ﯔ�C��P�}P{g�D옗@2�A�!7�P��sప�����m)Siex�4�� 4S�ԥ�@�0�*_��!��9�OmH��E�м�����妉�C,��5fⳡWz}���"�����I~�e�̟��BR�������Sj{o��qݹB*0��}N��ޙᶪ?P$j�Zּd�����=�P�=x�X��(6��I�q&���	��N��;3&�j��h�6��5��?DX4� {Nt`@`���M���^_ 5��J�i�"����HLC&��Y��6���1��BG��$��8Pj]��s�WaI.�#2�>s����� /�jl^�R$�F�cm�@P�CDk�U�"�A�8�~��fhMR2v���y��L�%.5���\ě~�B��䧜q��4^���k���-r*����R����\/���~��_xÐy{D;�sA���z-��-�= <�U�,�M:�X�ZU?i�� ��<�=S��'(�GdZt��\���iL1M���;�;���1��ܮA�x����t�%��b>?ӌbF���.����.O��]������X�z�\6~{c�)@�ɳ��+e��SE���򥣅/@��FK��v֫ڮ}+����i�J�Y�e�P�R)�c����q�Ct~����Hs>��G�d��LU�3�B�G������k���*�q{=���BV��A��'��`�������;��&�X6.G�j��}R)����al����C��q 43�hWȚp�Q[)�h/A	��6�~�'�Y+e�]�������HɒkX�3�ʙ/�OM�wV>���R�%,�x
�7��r�i6%D�!M@3L-m��]�W�b 3>��x�칩c_�Gшn*��`F1<���!9 ,K���Y��)���E�N�gVz̼�B�Yg\Kj�J�h�(�q�O��UX?��T����<`����y�@=u�6A����Ip�8�Vnp��C�����H%�Jx�rѻo��`��*��D�����5�+��7i<�Pѽ2��;]��������?���G��O���W������:�����S�-hvo��ck\ps���O��z��M�š�LHxAO?�f͍بs�A͎O�CIe`0�;`}�nYc��b���[�-�^1Y����E���q�X�޲^9`���	|�u���+V�J-5��w#�q,U���_�[�|������fHص���i�R�j ���#c:�к������p�q���8��g#0�C�gձ��! ��K��@�Q�x��D�����CɭG�DX���;
�t�9�=��MM.�Z�� <o��%a�6Y���%�vo��k�ު�Q�S~'a>��q:.��{����i���w��q5u�./.�A�"k��,Cbԣ�r�e�A(���/g����d�X����[��=*� ���j�ůa��{m>�$�##��_Kv���5]�!W�L�S�ы5e�����?LC�aޭ6Ts�G��d)�����������_���5Q�"�7 �<���V*2/Q��+�ͨ��A^~A�r�7��@�G��tVc�.���֓��$� u`	�����8����� ��dj�+���ѝ=?K9���hj��.-��9��>�Թ%�z��$�`�SjG{V7D.&��4)_�f%���x;���¬%>S�`[,�0��]Nљ��Z���9�����kT���1Ȋ+60ӌ��i��=��5���L�\j!�#2�l���a�}}6D�݁h��UQ���ya��cmЀ����l��qP&�T!��i)��M7j)g%bZ�	 ��^h�!J�/��(��pVȝXS�#Hב��1�S������|�	� �W�ZlL�Nn�P���b�=�3��m��ʃ"�#'�]�ŀ;�lv)����z��U���=�R�ή#�f��u�)Y��U �&�%o�u�!��E�Z@���m{M&l��!hu����T*�!�xon5T�j�P��-�t�CP��'O��؊�����\����%�n��&�����LQ<KSD;��Us��r-����?��A�� ��q�37ƭL��6;��m҂8��'�G,W��#��!2?���q�8ONJp���Hn��oH��� ���u]�a�����r����&"�+R�  OP1�n_��X��.���p�W� w�G�ت�Z�C���國��D�1�:�T��OĖ��YFL^��F��P�¼c[��ͻ���驞�o������i�"2쐼��>l�ӈL'��Et���[�I�,��x&���Kl�Mx���O����!.55��t4!����.YR���y��W]8[ל9�d,H���,�T��d�P�yW9[ntR�H����4&�
����Mj�T��+>O�s�� ����!"t��1�e.�����P6��U2hdJ���h h
$;�I�q�6�@U ���+��R]2`�uw��`	3�@A�/!��'?��e-�S��i�`���oX�f��6>Nǝ]�<s5s�K�*��U9s�]���n��$n���f��%�qN��Z�W�V�T���z$�v4��k�kg�i7��vV�D�:%Җ��f�:�B@޶�׊�zV
qd�~��o����Z$��}||w������.��	vG|�Q�� �(1 _M�N��1�8T�5�`�e<�����`M�6�)�,�AB�����z	q���i0�L���@sҀ�b�CO�;�h�!�F���`?u��/�ox�����IyWt��	�e�ɧ�K�Iy],� P01x��)0FQ�:NS��poזA�dI���ET�T��~%ٞ�|x��������<̟��c<�(5z�Ip��`��x`�/���d3��X�����rN��@�D�7��H���ǔs�rW̉�?���?79��N}���c���8��޲�j��Y���z��������\�k���l�0�z����,b+�N���i��,n��b )�N��k8f����ˌ���9P��
�'O,�
0!���QZ5�!���-g�,=Vj	��b���< a8�Qa��B��Ju]�G�Cd.���}o�-�bk�C_�J�!}�����(sڃD}�zJ
��-XfH�I�<LK�,U�_��-Mzp����O�hv�A�N ��r�ݤ�����n%�[s�D ܯP�:��22�(�����d
�uy8��K_y]�ֆ�j�Q�k~��Ҙ(��C=w�f-��?V�ΆUr�o��+��(fQW����̹KFA�/i��;����{��V4~?��Dh�%L���mc)����>Gd� ��������I�#%ï/�c�#�d<�Ğg0�ƺlɣ�U4^��$+X)K��s���2`���>Ƴ�A�.ߨ�>���Ppx[�
VFDӋ�_O]�r�0��pR	u�:�6rծ�үמ!���-�l�/���fM^is$.Ϫ$ʼ��=��7Ahͺ��ti��<���˒#C$#�{8��M�\Ff�nc:�\Yn�h��9]�������{���P�3�`�5n������9����e�m}�yc�GQ_8ו9��5G�Tsz�cɧ9�/��pU�}0lL�lc��'�� NВ(Z�r�"��g ��Ac
��ǞD6�����������^i!�Q���:�h�7��q��� ���,�0 P43�L��3[��z�Q�G�����:r��3��dU!��1����9�1�ȶiV&�>E۠L���l��i�E}�58���A���'S���E=�)(���-"�G��z�.+D�^��`=m�ϑ;��z�ɨ�;ҹ�N��M�������rPg�P�	���g��A^w���1�`��i0,�:���~i�R�7����oc�q����@"X��P�������y(��5�i���e��CX5Wwl�	5������#�.U�kP_�|e�<��Y��n�:���A���M�oٵ�l����R۞�,�����T���b��Č�6/�O�*��.@�b9T���/�Xtq	��m�E���b����Q�E��|�.*����1��@R�|����ehh�P��	����V���'�M��W���C�%uf���U��{z/��%�wxΡ(\���=�]EY��x��c�{}�3�}�h��+�L�g��+bOeM������C��]G=I�U�����'�V�B~ސ��$'G����
?pc	�8���])|�ױ[��\� B�\	��b��q�p�n�YP{NZPnuT�D��hi�{��WNȐ8�'�g,��9m�R�1F���u�Q�n㙀Ɣ��sU�AM�:�V[�㢇#���E����U-FDd�3���Q����1)���=��~�Ԙq(�%O�c�<�n��}cm�F��6V�s���eQz�MR��	ܓ�//@tH��(1�P,�}㖌#ә�(-�k0э[ MK�`ż����I1tu��P�%\�{6�ԬF�C��Ah@��ڎ�R3�x.��g��>�u� ���ޑ��Nh���C�55y�����hP�y��h:YE�o_᮪A��mG��B�o��x�M���~�
N��}��r�qhR>�|��?�n-@H2��f�h��D(�?oU[�X�5�8����ҕ4��R˩�v�lw����U���i���T!�"�� ������d�k-я�!y #f�.Dn�M`0^��@�:<�ożV{�
:���8_���˾n���<AB�>� �ׇ�p�o*8��u���A*E6��Ì~�O�M��y;�I"Գ ���8��V����=��F}���Z_I-�*r4�S䏐bqJ�l�V.i�X#����N�{�Ī�β��7ڊX�B���1YєUS�I\�8A��<+�ߺ÷����a�8-�2����2�~��~�6�>�̞�.2����5.��2{1(";�jӶ����0\��� �J�|���2FSz�'7F�w���~�hw���5���S[�?s�j���5�h�<�W�b�[���GY_�J[�'G.��?�o:�K
�z龜0�Z��L�=S�k�d�ǅ�&�)5{�Q������g*1%���zc.07Bs�-xm�%d�tv_��B��z������8D��?��Z�.����k%2P�ئs�fs��u'���|׃��W0kО̠ɓ��-C�ߌ�]�iZff(u��s���� V���p��6�����gگ- �к&]_N*��r&�I尰��1H/u#es*s��*L��Q��_��@H�)mrUHAp��ޞ����@�#��P�b]�f�z��X��\��\�)���ڻ[*k��W��|��i:��-�A�s��z���6wY	m��&�`�	�H�Y��˕�f����!$L��zi1j�` r�"$�6L���t�JJ�pKʀ�#*���y	ܾ)�e���G������r����i��u\3?0齐
Z}��x���~���g@��#�#|�Hl�:� {��6�E��}fi�+qļ����]t$ <Z,��9G*W?9�|�A���%^D�{�S;AR&-���������Us�"�Z�a��"�5�����dV�V%�4u��n�:�p�aTAm�^�1|�Bc;cz� ���s�8�P�z"iO�ݬ7���xV�x�z�(s� �]����N��Q��e0���-���yP�F]��B�1	���C2)�7���9`Ɖ&���,�N'ƹ��6|os_�?^�xrd�ܯNB�[���&γ-j����tsۧq�L ���8O�����yz�����It�ع�`p��?��*��8��)��W*tb�:ƾ^M�E@�W)�9�&٧)��`f|��pzqc�*�T�(���ĝ�"kL�>���1��|$ӕ���*�����6��u�J,_u�,l�[�V�[��3�4Dx0��vMf;g��uL�hrI90](4`��+}���c��QK%����V1��3ŏ�C��i,	s��߱������~e]�)˸�Be�]BL��&1C�E�>�}&�6S�Y|p�-����S;}u��CU$��AȤ��V�fã);Ob6�رb���&��ti���=������M<�҄%<)�����o+p�7��Z^��N:�_i'�|��~�YS7in�5��gt>9X-��
�%d%�Jf	��S7���_͊Y^�)�Id+����m��ǎN�eR7��k�vr�ksc��G~3	.�4�w�&���h�C�,���<�W��Z�*��dx/�m.��Hg�d�܇��#���خT�8�tg�q��9iU
��`�����;_ٛ�Y�1Jc<��{��?k�b� �іَ�lCD W��/�R�AL�}3�)dj�A��lS���m�i��\�R��b�w��{����k���.+�J���5e��l�#;�F�����R��!��g���uhzY��'�I���ar�@Q�9�
�V��ʙ�>P���I���jR�/�H�<�s�l+����=�+L7R�w�&gH��� �\ǱM�݃�����8�b	��k|�g��״F�c���:*�˾z7%���p�.��U�.���7-�7zcvd�`���� t�[kZ
�/mX���>M��t���&,�jq��֧ �LIh�2�&�}����o������-�|�vǫ
��_aeўʸdY�h�=�v9��W��9�� �_
��w;����^d*<Y.>�Q
e�O��΁���3�f�,��=X,��]#���%&x)ߵn�dK6���;ZH?(u��gNG狉X$ń�.�1wӘ*z0h�.ӕc{y�i��2�΃;-a,8r0��<2g7��l&���0�F{A��q���-�{�p2�r'k�/]Z�L��Fx���6̺ *�<������7 �5C�����2�����i�"(�:f�}֮��C0��뺭4p:�^��D���瀕�:r���A��T<�r�/�C��b��99-�87���b�Y�V����ȀD7�W�7*�FQ��y���ym��r�妙�B���	<��ۻ�zg�VI���-,�tr��|�[�������.�e%���Đ��E�R7�/\O��ol��1C��c���(����Y�$"*�tL�7��R��;�o~	��/��F��9t�c	.���ԟBŃ/y!9!�ߑف:0�$�e�b��rP��܅J�� 
�.z���T�DÓ_͓�k��Q��؉֓Р'��8��ݎ�g���)l "�;|��E���fyw!��j x�$�V�J�����5�h�*�;�w�@% ���ai�a����yX��LX}�Aq�,q���Z�8�&�!3��x40���{�ˋ�*��d�F�����g�ς�&����
�Ҽ�k/r��,��i�%8�t�QB�:�o�|�m|���|ܺ�z�q��M�C�D Z�sW#ٸd�g�-�	�l�d�1�����D�ќ[��r=eV���Y��q�F�_��e��"�흛yP	Uw�)0,ov��V�y��"5?U�>�}_q��py�U�4HT_��QD[ˈ/|�M�����1��+.`��B�/��%V��ga����L��Fc�yh�V1�O�D	~`z��h����Uňm����i�<x�C��@�>���n���Pd@$�\��)��6��Z��U����a�a�9~j�i��:�'�X��HU�FD6���1ɍ	}�5�h�b@��}���Gp�"�Cy��T�%��І��GU��\8��;N%�*�A�� c&P�
�Mp���ހ��K�hqx�{n�]F�����_U1B�[3궾��U�
+{��SJ|�TX��h�0(�ĕi}��{ ��ɏ���% g��:NF���<�@��$~!0���}>�s���V��+�s�N�$)�;�W�V.��$6��=�0M N�D�T&g����"��*����5p�0x����nb�o����E�O=���E����s��~�9�'�L���%=�q����$R�Q�::q�1����p�[>��/�*5������/��o� �����m�#�΀�],&,z7[��^}��Y�t)�{F���b��n�hw�:�e42�ӵ���X���0�TG�U�m�H�F�w ��.M'���A���ďׇ��?����z�넔�H)}��+5=�*~��,6��u Y���>���Ix�����N}\�:9V��c��?����җ���^�9	"��"��H�K���"���D�j셕���D[����i>yѤ��T� 'p�Ć#]@�j܏�i�>��C���M*D�(Q�`�F�[��S/N0����FB_����!Hh�b�I�n��&1}��P5T)B֞�"bvx-�~���CNz����"Y�q���E���_���0����?a�3��Ө��+�b�0GJ�aN:���t��Y�t���RIG)�i]��ȴ�論�����i��J��`К��eCr���玧5eEa��`�^8�G��N�1�'��3JT��*r��O�ΎGsv���V�K�J$�
�����`Pk0z�
��≠��I�@���e��BZ�o���E�>X�N��A�q�L��@d�т�U�V��EPN�A��j�ο�
"I���>�yF���T�6^ٺڣ���d-.bW�����hѨ�Z���up������]'ly�����0k^�U�j�3��Bv����ǖ��JG�$�ӻ)�������*.�����	�ox�D����x]4���jj�%m�~Q�zϼ ]�����U�pRl����K	��fwgeje�_\���C�(����Jcj��[�P{��۹�ٔ1A?��4-���a��K�^���A��)O�͞�GgG�`ο�����=��8��Mu�=��e�1� ���5����-�'@"C��x�ۋ5�.�u�iNl���
�0��T���Z��[lT�X�4����K�4�\pɀ���/T��=��#��t���l=l+��-��^�O�wD�>��R�OP��7��JC�k�Hg��A�U4z����EZ҉KF�?(����EUV��5�[ 3f����Џa�/H�� �BьXΐ=^�B�;�P!��VYK�מDX��U,_����pX�[�9��_ZZ�h��7a-c���c�ֺ�9fn���u)P5�b#�t�=�XY��ëY����{�-�1�;R�C�A`����!Y������(qu��� #F�6/��Uݦ��ωGW2x��5dW��={�\��h�B��te��w�q���д�Ӵ(�d��L�A�9��HT:�^�}�`{B%!��8GA��rBB�p�X�c��]�{׍������4�gV
F-�iX?����wt�7��$v�fꄃsU��؈�y��rSWmi�Im,bV�Io�* =6�rKO�w�c�"�j��	�7�mߥ�`h����30�o�Y���
]�Ώ���.�2��i�4Vk.x��(.�]az�#������庩��Kk�t�e^��z��L�ߚq��?�{E�.ޏ	�2���|�� ��Y�3���Ȁ#U'�����/�����V�~�z�M�ťl�L��\�Mt���
@�|U�Z�@t#9��-rئX&�6Ifɷd�˥O��s�������t���}�eB�Rhx� �|�fX����j�ޡD-���ZST�����F������ﷱ�5����9�9(��I_҈�� |m�*%؇���sm��S��X����u�C˺�U���r��2�/�����������F�Л��G��e�Q��Wf��阪��wZ0��D��C%�!����_�w�:PΤ!,S�����7��3���0�=����w�X�J_덣!5�Ev_5��z^�"�~k4 ��)g�?y�4��%aW��_�U����B�5������hCi�^��[��c�٤�Ԝ�A�
��>l`Y8^�?}���*��[f�����+C97�v�����ړ�?�CK�\E��u��i8<9;�.�.�;!Y$��Ȃ�>I.�J��AZAP|��u�pH. ��0�nBLG�[/FK4��к�4�h��{#��������.�7�?�f�8�̧�ۧa���u�FY\���i���ɭJ}����O-6��z����� 0�g�*2�칭%^��{��e&c���0�ҿֵk�v���[U�*���eV�N< E~.� ��+�8�S��h�wp��ؕ*��]�p�َ�0�%�P��d�F��k�X��)�c�U���yP�`":��� ��j��ݓ�,{Q��%�&2q
>��������"��%"��V��!�A4�t�7��μ�ܓ��'���D�~��;��TF
��piI�u�� '�����S���}$���UB��Ф���d�m���q�L��)9��Xsl�T,?t�.94�IB�3o��P�+4g�j�/���r��G���0_7��wY�ա@b��%t�#�Tx�Eu�����^gx>=�!�)���gr �6dV�R^�b�n�x�]G�̦�1��c\:"��}c'�'�Z��a��d��}���s~rxǵ9������nӓ����v<J���`"�ɰ�h�����R[[���(�y�y�:>F��N�!=���MC��F@T����ҿ�[.���\|�\��"p{a��Ԇ���~9S,
љ�֠g���/�=� _�;�P��ֶ�ƀm|C����+�����~��P����2 !�U�L��ڪ��zTe?�;�//��)N��*fT�"5�y¨S�Q���>��0����%Yƶ^� �/Vh����ﭓ�Lf��|�1��D�`�׸�=���w�ˈ�8#���4
OgI��y�[�?�m��D崿cTi�~��;g=���
Y�7"Ü}��w,���"�j���G�4 ��E�w���RO5c�4J_����?����މ�T������W���_q��"c�	1h�N5���  �t���Pi ���%x����<����l!�:D� �]�����0��ǟ�˽�5��-*sx�f��-A/AR�dQZ�\vI�O��.^��^VoѠ�.G	�X �j>y9-���6�e�Y=�i�OYl� �
�^^��U��3m=:f�`�#�4�mQt6�u���ϣ�qV�v�L�*o���wR5#���ϐ|2��׉qIK{C4�뜫�{�EW!���>g���b�I������Pd���?�
vL$�qQ���a�y���uҳ	�W���' ���m���H�����!�}&F�S }0z�Vo����sG�@(π;�u��D'��U�E�Ʋ�xBu�f�U%�8ՔQ�i���Puɜ 8��*o=�U�i�d��%�f��-;�_�'��8���i����۲Q�;_��-Z��2KPȦV,��.����X�:qE��~Ӳ�+P`=i�R��薪<�S����}c\}�~�����'����Ends�IrUn���[o䞊�U"�c�<�W�Ur�4s���@"㯟F�1`G�6$p����Z�/�	(���,���ؘ�|[�bU�<���@��ߣ��#�	0���؊~t�KXU5j@��W�ı��k)1�{����~�P�H�HwלL���w���6�!�Fh@x�+F���C)~}�]r�^%�*!���h���4WXSІ1t*[G�Z��\Z�fȏ�ɷDub)P�P<��&����(1E�?"ȴ`8�`�(Q)�1����
_����q�ϼ8���}C��#IɃ����[����T<<�d����*�/���s��f�o�'!���s��k��(Q�w;$�\񹲩	�71�I��d��{���3B��9b��y��UkH�^v=
l�����e݆�D���1��b5�����?;��#��.��nTg!��7��M�*����Q���*șjr��o��݂8HFw�ȧ-�`�|Y�;�N�q�s�D`��k#��W���W�*a֔+�فR�?��ߴ��π���K���e��3c�N�<�-��F�+`�m�t5`ȱ!39�П���oY��iSz��O�o�K�ε�}�z�0���d����X�_���4>d�'ƅn\���(x���Cb��W
����`��Z���_eZӓ���������Vj��4�ɬ{<�ŕ��7%�e�x5&߷V�T>�C��Ⱦ"�;c)rͧ�ilOҘ�Öj�]����M{wm���{�O�Z8�ch��9�@!)���?Lـs�uW�`��-8|fU�et =߂1��VP�|���O�A�`�]�x�1*�T'�G u�Rb�
>�`YA�vj������;�\�j43s6Z�j�8|���K���(���l1��$4&��X��f��1�,�>�(�ssA<�o=v��c��5�+0���H�l����;
Cz*>��X|)�����%�Ъ�-���?-'�Ux1�6v�l֠ _Ȍ�����Zv��G>��rM��M���G͈������H�-O�������R��} ��s�[��>KH�6�S:NO���U��~�g�u@�#�)Tn8��#���ˠ�<�ԖT�53����g<��0"��n'k��,R\ o]����a�U;@Ι��An�[7Ǽ��"��Wuk-���_ w鮛��%�	0�>�|a���>�ˏB�v*���w�Z#�v��R�l�k	b�;�//]��_n='<�iy�Ջ�t����JW&�Z	��,�z���:�%�u��i�o|�U�8��D��y���z���X�8D$H�}�͋�+��{	��i�`����)y<ph��ڵ��s4��YF�Dջ�h����%�ǝ��	��J�e6?l�4� (F��2xL<�Mp��2��3T+UFm�(oow[��m1�2�2z[6A����GIb=��fi�p[1pL�ν�f��l]*D� w�&ui�Ob��uu����͝�o�պ����Z��H=>*�(�5H>�^�v5yH�^�4���p��t]�ig95�1�H�]�k���_�NF���H��>�rQ�C������wI���&ZyUո�r&C��U��i�"�U��.�p�*�8�|H+�W�(E��R��U���	��V!�d�R�����:
כl6��Yg<`�t����x�����1zU۲+\��V<��[�>E�3L:�B%�h9W��'��?P�L�ȏ^�y7<�-s�^n�7���*�"����Ou����?�����e.�mo�7*	bߞ��W&V/���������9��:A���B�B>�M>��O�)����V�BĘG���4���C�lmk����K�Y�OH�+/��<|G�L}T����_���e����Ci�����$@�����Ő+���������7����d+�"���oS���)ܞ�w��9��ƨ�I5:�]E����q����w֤��^�׳ػt�ɒc)�mRw�������/BH=3�Ρ6c���n����Q�}���1r��r�X���Oɭ�BM_�M9ϻ�<�{L���x��`6N���[�,��ZsL����I(��	�zu>)�6z2��@a	���T��F��'���Y����eȝ�>g� 2W*η��K���7{y�A�XsR.�>%��Nd�*�Z�t��6���Á�f��&�|��yl�<M��R�5��L�tP�l�=�Gh�#z����ꮯ���c͙��>��
�����O{���+��n��(�88�I�r��@����=�`����۸,�Aʽ��V�èG�C@�(w�G��~�)�*��y���4L)�q���/S�L��g�q7���*!��XЊ��E"hSӏk-�� ,-��6�>�̰�'�M@���&��C��eV_RM�������]TB��:2�ט?$y��a�Z��)M+s�mk�)}8�-������W��-�����M�	5z���g:�Rr뙀���'�F\�	�3��,�R�7b����Z��&(���*�#�d�� �z��R�
v�@r��rEm�Sb�)bW��g��rz��l"Gk��@��1��=�v¼�R��"AB\�r�QH���-n>�TK�ܢ�����e#��N�K��j�O�]��=�S�Ғ����:rhPy������u]|��Dح:������S�3Ή��O����7�ۗ^`/�Jq��Pn9�Q/O�@���K�;�1S���&~�3�T���4f�^�������W���RJ_��Ō�f�4w.8#G#_}(D���/O����T�#����z:�Z�L��'֬���Ld�v�nlF�:L^���4���N�T��Z֬���`-�C���ײ���Ķ��^s?� co�H�����V�¯@��2Ο/�YL��0���a%O�ORX#�-�W��{�N�����Ƣ
�v�Ʌ��rjlK�VP�<�qaafz�=�M��n�����;������6]	?����M�|Np�]�z�G\�&��`�>�xT�D���/�uho���*�6A�~-zO��[���Y4�(��T���Y,X�7Bn��?[=�ϔ�+:���8^<�z.n��2]{�3�m .�j�ib��B�Hs5�Ȧ��g7|wa���u��b��f��a(�S�0�O���cELdz�|���#13������i��@Uk��-r{A����T��d�X_J3�>g��38�/�<����S��=5l��(���x(���cǸ�S�uP�!�����`d�з�s�M⌡P��O��^������u�nٞ$�O���־g2l���$�)���}c��/7Ѓ#$ѧ��g���������cR�t3&�Ae�u�L�b�@�;��8�.V'�~��1���i<]`^#�4��m�����ns�u]}�O�6��A���m�qh�ك�����k�A;�ȥ���O~��AD���+�@>��<gU��^�o��҉I٢���H(�0��n���G���g9 0�����|�  �RxS��Ϥrr{�1Q4�m���hVex5��b�0AL���U���ڀ�^�F�@�$�@@&~��\X�}�����Tތ��џ5������20� h�V#��[d�����"�ϝ(�Tˢ�3Y�p?	̙������Jeǐ���8ڧC�����<B�8]4'Y�3g�j���0���O� ��׮���oܺş��R�Ў�W����ˡC6������Q��?M�tՃ���޾��Vw����"��v�]�i,���ʖd?��P��C�b��~�@�=�X3B� oFI5Z�A�6QÑ�-~��uʭ�rս�qӃ�����@k��ػ��1]���ɀd6��	��5.7~h+�=�@eZ�Z��?O�M"�sp����M�oL��WB�+g�:cg��G�!��[��s�ߨ�1�����W��(t}��O��V�w�O��1��#UjeH��_�0�M�D���ɎGr�2�m�/����@/l�@��dK�!o��x���߄�Ԇ	��i7p��~�)���.��T')Z��}R�2��Ȇn�F�i9����LZ�&f��4#F�]�O�?B��ە(���nw2?���wU�o���b*d�sB���ۗbm���0+��蜀*��֭q~��HXj�C�q���2���]Y��Pu$:z��A�:�p8G=����=oA3���x}��K��@ʽ�xɅ��IW!�cp	��-�L���̬���D��'�!�F��Am��6|�?��*�����cZ:b]�,��Vi�{w���
k�&N�2����	������� c,��`�?'�w����~�-�p�"u@,D��د�o�E�ܷ1F�T���/s���۔��xb�z��,�>ی7IN��d�"\�#Dd����% '�[$C|��ν.������
���@4;���)�֚���$03����z�9�=�ͲK����UlgÍ���rܬ���&�%q��q�Ǭ��"f0`<)��f4cu���U�ư'��f��6 L��{�wm�
Ѭ����@�R~�|��VԢJ����CYa'`\t��чh���䌭햮��I��y��lM�'�����6l�}�I0��ׁK_Y�.u�əV�7�6̋���5yΆ��l�
	����rZ6S�A��t����l�:eϾc��6Ԑ�7��Gf.�h����ժ M�����6g���M�q$gW9� �~8}j@)X�
I/S�e��$��)���.��C<�	;<z��oU�Z6��^�aq���l�l�O�hJ/�M�I8:��&��4ËDf���d�U��
m1��E%X��b�	Ѝ��F��B��I���Ge�;�m}��KU�Y\��Ew��3b�g�2�m����G~�T��iW�Iv�79�r�I`��o���ڙ�K�!?�����~e�kRe�����g�}"��ⷖc8=�~TIU�_W��8poOY�?��d��n���ܟ�֬��_����ސf"��81���fvв��&(�Sӑ�2�,�O5P[�!�h�Q`
l�T�=4qI��"M���!��Oh?�c<�)�z=�����J P5U^�>�n!��0�'�o�wk� �I3��DBR��6:vkܼo�����ٹ�?��R�s�f�(V=��Z�o�DN�:φ��&1�DX]���b��$t(4B�S�W�����FU�+^t��ފ9Z�s��m9
�ךr�?�8p�~8@�TT�(\0�U��7��S"�8�@g
$q ��{�z�c{z��-Ȑ��k	�VPžf<o�żǇi���oǾנ�EA'��M	�� ���r�6m$F*��_�`��(IEL�ۡ��(-��S���Lg.=Q�T�ׂ�(���;�N��V��t���b��{�ďo�~�f���	~L�V��c*�XDS���7U�,�S����������u�~Q,�._�>we�C�R'сH)��7�
%mOS��*dK��������_RqeO�fs7D�+�B�\Z�M#5
��oE�Hw%W��GC=7�����"$l4��$��\�������ˑM���W���N�!::��Ռn���$�q�������*곌x�,�>�X�ͺք�Ox�3St���	���e
�ucg�۬�yɐ7Y���P#g)�H�cBgd�c9��I�r#?��9��l�g�i�iW�3ud�ߏ?z*j}��� ����P�N/�F;��SHmv���4Z�׾-������q�\$��T�q��b��(�X����cQh1d*y��I�<�{����S.:qKFF�W
Ys+h�^U#r�VX�ɣQ�t5Y�6��q��}iJ����g�^���Zcp�-��S��.�9�"k������)'�&�b�"�O+
\j�nG��Q9��pu����^q4�8w|�����(�:�l{&�c����{��f����MG�խ(�j>8���)GM��<i�� ا��g�����@{�̙$S+��rfS�Crdm�Ά�-���`�2�6`y쭅���Ѕюuc�v��� �˽g����.9>-,c]����!L�&�cf����o+�U-��HM�>⹲�"�`�	�)��H|؄���쇊��Ê�;2������턌��~D�V�E�l3^���iA�#Q�8җ2X�a^F�MA�Z),��Z,�`{(I+�y^��шr2*#�{<Ո8�FN1Pp�xv��ej��&5�	ޱ�t¯4�JO�Q<$ɔkI��M	%��Ms���9� �$RA�ѹ��fG���; �?�R%�If1��w:_����W;����h1g�ӯDkM'ނ�BP��~m��5K��`jǼ�I���dL��YJC�Ӏ竪��oמ���vì�FDh�Ҥ�c�n77���$��4orz,��J�Mo��1 �5�k���L	�j�����=��Q����t��a��X;�@�>��)j�z��O�To���(`���|��fz1Ż7&�����F��.v����o��w)K���L�EM�D4�Qcq���.]!��#�~�X��ydC���r1��6�9*�r���#�xa5��+y��vRPc���Y�N]��B�������U�@��sF�mK�,*��`#p \��ۿ-i��*!;�vl ��n!�E��:�;����z��]DY��]��=�Ϙ�P��C�Z[;���c懘�*o.Qf0 ^И2���^�i?��d�!���v�D�g��&�; Z C+g�g��!@	�d4��+����q����^`O�H0�[�ei�fO��f��������	b/��%D�:*��v�źy%A���"��W��Z�:5>	��\0FM�7V�~�%Z�=����k�g���Q��`7�7X�B��ۨ��r��\g�Cz},��*+�������ʝ΋znwlbʔ��'B��C�����|~L��ui�p�a@:{�/ ��F&��xtj�*���r���$F��̋���A�&�Z:�| aP�(CC.l�vd������6�j	��z�&ԋfuŞ���5J�����M�Q#i1.xr$����WF�:��JXcD�+���YfHy��E����Uj$A5�X�$�	��D�1�?��fY1îSf��"�Z'<"��G�_�Z��<C%h�y��((�|�����`�A���zA�Y
j��@���bXF^�+��ܰT�&���p���4Z���(�D�L�B��f��[� s�v*8Pxy���o��C��h�z*�8x��ܾ5��;��J���g��_�!�י�K��E����-�1�`U6�+j�������x�<�2�&��o�"�؝�%����>��P�@�j����0��z8��C~9l�M�%n���ֲ�/��POPd�z�|�x���l	���D��յ�<��˓l���׫&k�3� �A���x����mB�T�\����n#fߴ�C����.W�#Q{:����#7]��9�H�)h�ҮK�iQ��X�}˧��'j�h�^��	���_���h]�1ZN�g��&�W$�좷k�``;��4J@k�V�Q1gSUh}��'p�`D�'oI� �8#�Jl���\��_3=+�OB��er:��W��*�[y��W�l
��[�Y��,�>V�s��:�E�r�������_ɛ������@��S�r�-Qw��]y �����׆��5,%�d�2��C3r�;�FA��m4�bS_�s�� �%A!t����@ItԌ*�}8�@��
Q�^�O�CeI��:�^��~o�k���qi�)�����d�G k�d���@[1eaE{	_�D�!��(_a�c���a�s���m5��o'J0�,�����qޛ��^���hvT9��EQb��d~��/M���|�7e���ХNq�x�9�z5� ���b��>�
Dw[~p~�Y-�\��YUG��T�.����M��vCj0�<>r�^B�W��6�5!(b�ǊW����ɘj�e᮳|0�Y{���Fz�����'���W匵�y��`4�� �⒑���ą4s�L ��X��'jw�7��hg�!s�Ki�3��V�X������<�o|�_���x�V��LhZ��$}�H�H��8�
�$���i��6e;
(����%�#R[�WV�nI���X#��?��Èoz*LT_��<�'$�� ��5�V�FͰ�-�v��r�O+7��G���d�e��V,��$]!�(II��\B�����J2B�kIk���7�S"�|������&p����	:�^�B��Cܼ,�|��]|^�}�!��Tش��)!"�L/��r��GM�k�R�׾4�]�iv�A�����d)E�C �ç�����Ug���pr��T��o~����NP%4D�ä��&}���̲�8�Q:�0,r0�p9�E���0�h�k6���;[�]>���ѥ!�-[zoo�e������Jg?
��r������qų��/3#��	?QŶ������ͼQ�����d��i����m.+jRp(`>n�MM�``aO}��I�{��h���M~"d��6�ʄ/�(6Ps�d�6�A�����������6��[٧j����m���X��Rم�>�UYް���q�~ц��Yxa� #(����!;2�:P�A�1)w���ĳ�Duҥ �6C�R_��.��������`�zd��EU/��3q�%(Ş��h-���nӷ8Ket�A�h9aFm�<���u��R�Î�P_��"S���r�&�0}	���Ԑ0E�������f]�j�6�0]���
2��&��I�����q����J�w'�8�Q:�u49V%?�]ęôُ�#��j�*�T�����Y��9�k�cZ�����ȗ81����XQ�Z��kd�R�������E
(<���NNp����i�7�=�I'����̍j^QU;kM��Ę,���?�^G+=��#7������[�cq3�i[:���G�x���ep��h�p����N{�Nѯď����-L���
>�ӌ�=)�Ē],o��:�J�/�<Q{��}r�K.r�֦�(!nO�sU��bG������x�OI�"t��t��a�FRșP�����2��.NWܪ��'p�;$p����A������w+iH�2�-W������Ǔ���=�����x� /��`��&��x��f����P��σ�����nR�r�Խ�V0�f�^��Du��h�#����A����J��`2�K �Zh�0,��H b����Z�$��C��8��^�|8Vџ	�
V��o>����2��vCN�vcS��*�w�����g�fb�4�l���9&o6�F�S�R��B����zo�O#�H%�����=�Ǩ�X�<���y�z���!3�'��1*��P�1�~��)��X����a����#e��\�� �zhT���C̰Tכ:na�x����}F��B�C�hkӍ�嘽��p�1�r �ףѧtĎ�ȝk
��!gcs�L)�
\�u#������r ��k��[��i%7K�n�:��Ⱦ��c��97�A0w��3�?���7�un-�J�gf�^D�y3B�@��^�����TFl���q�~�ϳ�u�M���N=<-����t+̹p-� Y���F6]�D�!J��o�0eu{@Xi|�7w#3���N��H��߂:�#���N��`Kgm��=�؊PN�-��\�����eAѥ�-]�bz��j�L{"yN�K)�x^Y_���
̌�չ��4�Ro� �E��1�Y)�	�N7���4��?�!�ȶ�Q�2���a�(��o���r1������YQ</._F��U� �Or���ɫ���#�/�����1�m:/�צ��{ X����>h��Z�e���}:�Zf�~+$f����a� _��O�|Jz+6���t[���φ��O���A ο����8CW�&L����1�c/Q�ף�ƾ�����q�f6\o ���W�T�~[黭J<W3�=�WVe�#qأB��t�~D�F���^�6�+3l�-Y���Ya�U��V�~~o�v���*t��kݐ$Vm�Gy^�Ǒ��̊�{iV�tO�EQ�p&���`C,��҃̂t���Ӥ�r���G��2�yEGH�p����`���l�+J悳����!�"n�>��##CTc�2�v�}n�^�]T0�t���0���ƫ��C��Hdv�3������l8��v ���ό<
dok��U@�ߏ��v��Ĭ*�&TT��F��t�Mk�IE�7HP� q�~>�K�9�7ipB�#�a��2�
��cq�=J�sd���hX뼬7�@aPG�����f��|��J���q�dG�p�C��Ԕ����įw�woRջ�?��1G7��q�SnӢ޸W�M���u�����t �nq~�����6(�X���N��O߾ʏB fd�)�<^��
*���������R剰�=؋1 �˩$瘋����R)-����H�Q2�k@[�?�(��?Onm��\ԯY��"#�Cg�{�:���Q� Q��h������a�:� ��+�Y]'I��K��� ̀VOᮓ��c��̛���,�Q��J�#^e
�k�k��T�^��d�7�u�4$��}��T��g9bSY=��(tюX~s��1�nڥ.�����!4���pו^@{5�-��m�-y�7�UG-��h�ت�}r�m���C����u=���a�f���5�J�?kO��%�ez��J��4�+f"�q�i�R���L�͂*g� nԻ�.�)w
4�9�����[��d�����b�(�?�6^`�rN�OS�cD�YK�`~�9&׬>M�/Z�{��)�#�z(���;���!�����֝ԏ�ĽD�g� �ʄ�U�IƫL��oJ:�h,{�l���*��V|}" ��ԑ=KnD���!�?�@�`��;����u$�<�+�p��r�{�ܮ��BP���3j��B��HKX�����	U�LcJU�p1a��5(�X)M}m � 4.P���e˻�Du���n:�rz��i��_C_N+o��B�1���GX����(p�Ϋ%����!��6
ƺKE2���?"���s��o{��7���� 7�e�� ��h�$���L=� �08��S�H��O4z�'�v5
�K[���-���[��a�u�u�t��j�hHHE��2:8��Tv:{r:���\���rpM�M�#��b�����~�w����Fj�3u��d߶1�xRn���7�p^�#��԰�E�t)��@F�B��}�'�?���T({��x@���2؜uLT+46�:?���U�A������i�>������6ί,���z��85p����d{-��Zn�GW�u�~ecP��X�\#�-<���qn��9���༶�u%��>ȃO�O�>7K&���fQ4Vy�p���wEź�=.�c�B�A ��ؙ�5_01I � ��:S�e.�ɩ����+��4����GAG�uy$c�\NQl�"hP�W�����5�I&ܼN��Xs��z�pJ�SH|��:2�=7]{���̢Pe�m��]t�X��۠�2�K�I�50[���ǟ��\���m���JS�p�y�G��9h,ie_ʩQ����a8ΚN���BB�)h������\����Gu� MGc����9>�j`��#�-�$f�b^RC��J���:ӄJ;�Y����#��r���� �6��:6��[0g|IB��O��iR EXi�hR��B��k�����$Q���ypU��Ƣ�N=���	f��vf�B��)fc��?�k��5x�F�|��<�m���<����4��E-�#K?�}�������y�uB��\b���%�x�ۭp}*�몡
�� u/|P�3���1���{aN��O*�ݩ�߆��JH.8t�.�H��2e��w#
sI/9�QZ�Kf�Ț��R63v�>�a�x�(�soo XAl��YLNW����?^LҬ�� �$<Y)���X���]���ި���>2�~7���dM=��׶���]t-�C���oҨx�ur�T�H_�--p&P�{b��V�<oı6�f74X{���S�.R�;�\棣^�EyV-o����1Ȧ���5�Q��% �_�xx�r�]�S�"�cˈ~g%�\�b����v��u}���}��k(zZ�pVX|��A}� *�k��|ػ��'N��F��~�_.ow���f��A��`�tv۰0����Ekv��tʍ�����U?y?4]�5q�+ﬥ��D�<�WD�)�.��xm��G��TV+*��i�;�V�e;��>��e=�� ά��0p=9�I;6��>g׶��Se�!�}��>�#��c�Ajrk�3�9Y,��0�xHl����왻Pk���LF�]Y=M��^�qV1�Cj۸<�=��oe�Q�Dl�*�#�1�)�4�I�.����n�%����x-�����C�y�����5%�?�[�i�� F�����5	f�����
jW�ZR����q��гdҼ����m}��P]�{P�75�P��
���N��E�'�K"�I��$2&�S��'��?8���}LC����;Ջ���?���N#���J��������H���?�(�7:�f��$h�/���y!8���:����2�<�аQU�X����1��9ʝb����a��L�����嶒ӂ��N=\(�6����@�6���#ʉ���o����S�\�6~'	�!�oYq���JS�E�/�E�@ K
�N��u�:Sw�CKt�ގpi��8��|h9� ���ų�~�\�4������Yn���k�����H��$�]yX�?U�����/Lb&Pv�.O�+��uX7��y�A�n=�� ��#n�G?S��bi�u��s/{
��Z��(��9�5�1�f��ij;;7��A4�?�\T�GT��j(�������3�yc�"=_�4)�Ư�O�Fm������XX��Zm2
C�����Q#}��7��c֥i��9}ˣoZ��|Bw�<g���:93������� ���ʋ���;2֮����)s���Iy�׾��ex��N$f�ns�Pŏq�^�%Ӿ �i�Y
 �Lh�󕱓�b4}_"h�3��NgC�ѥ�PR��j��ub���,�n��3����i������`�G'���G�vև���m&>x{r�|c��ͼdT&~�b�O�ŭM��)nY��U�����������z=�G��Z�)K���]>���`(��n��ϕ��F�Cd&�x�C����ֳ��+]@s3��5e'�P������a�l���'#e��Qp�4vɰ�z��Dw���Cִ^t��V~�x���&tI�\��k>gx.���������,-�����^�t��bL����0Qn��~��fq�h3�`�T�y�~��^�O��|����m|Z�Q6u�����������U/�2!�Oa�grv�`�'�7!��ct��}�@H!��[�!�~7�O!EM��5�Eh�	`�p���>�p�]w�C��}����*%�bB!��]3 ���ó���Pw?�j]����n|�J���뮞��y��A`g!L�J��Y�\�|�f ~��&��D�+_���T_
`owK��=�pI�{�������X7��j|Q�Ӯ��[���P��Vc��`�ôq�>���7�C�����3�J.���p�lK�=��f�uAO����� 9FC��y�V����IL�8�n��4بG�_�+�??Q�B"R+�H���/E���k�>W扃�\���KI��f�ʮ�����5y�4�_��*x8�O�ޘ�߇{���A�vd^��o-����#|}R�l��(�"�> z�dg��"in��#��
56���o���Dx�PV(��˹V�Q����a��澀�Hk��ֱ���A��5}�$i��g���ç>D�\��2��h�	�N�v��Q8^��=kn��?�ۑa����Cm�y��po1�\��U𗍡
��vm~G�O:��'�a��<:�NA�"Y1]��d7��"���3Î����HD9W�5��䁝a�Ob񲮎���)�N�_hQ#^Y�0�M���BE*���9�2�F^���=I�"7��o�P~�'�ݒ�Kb�mRr���K����x9����^�
�y�|K݇��x�,of���Ę�Qq)�(D��R,���@���4�2��i��WC�W����v�͊����s�N�Gtq���n)C�O�Q.N%���Ġ.&a�=T38K�S5	�ǉ1�����Xb��7������"?F^N4ً�׺�]U
�q�9��7(��_#�V��@n(�ԏz� 6���=>����0���xH�G�q݉/�b��|-$��E�I������)������W>�g������2')�����%�m|Ə�+����O�?M9�:�`�e�=R���R����k��n�*��+��W�����8?+&X�<�a7�@5�Mj���U��ZYU�fv���ZMDw�)bD�U�aV�F�}l��Q�"��Y��t��7�M{���8��!Rc� m�l�@%<}�Â!��4����������%����0��"5R���`��G�v���f�VqA�}�V�?�ʨ@A������y[�տ0M7Q�cq4:�ן��>��Y5�~��bQW���)��HN��HȵG���e(��8����#3,�V�]��)��=�#�i 7�'E��[,��a����5zH�$���ű�� B�B����^����ş�
�����#��U]�3tb��>����N�	I�TA}�a�I�g/�6�F�ᝈ�.d�^𻕴P�]D�[��J�k�����n��v�v�t7"��(y�$�L*D��I��.�k�AֲPEu����.�)"�� n��1��m���o���gH�7�ޯY���o�܁�I��	ҟY�'�y���c�$�>�Vr*�n9_����x�!�hɝ�\YU� �&���Um&_9�s�*)�����o������<D���䰜1u��:duR]���h�=�W5��8�/^P�8�ߒ( �c-�S�Ι�B�ݨ3R�r�Q�"^�jށ��]��״����5���n/������u)�v������t�ܲ"7?.qhU'"�}u!�L��u�Id7&8/�+�X��"����y�4��gr���`�m~���+H�)!�)��S,͑��=߰��L��<]X;�e�1umq#�k��IR����i�2���(�ݖ�ٕ�\���\}�	��<w[���5R=�w�`��qY4��M*��h(α%k-�Ul�����������j�ɝ� �꽊�U��5��{CM*��^��m
(��N���㰳�:�:)Z�}uړ])���Op�+$Z��$�FI�6V��B2'e�i�ϲ>�:%���%;�� ���(�@���R�gQ"��l����)�E��g.��X�*�&��>�t����l֖�
��ztǇT��Y0 ��p[�o	�d�#���:>��/�9�2nڈ�(�sF�/�'̔-O�<�rbK���<+�F%'������"]�WU�/.�aȱG��(Ɖ��2�ݥ_T-���!�\�+շ$����D�"aI�^�ˊj�qe����`�d���f��l�����uZ�o��i�az�4rm�LT��e�⠂������6���d�`$�����U~���f8�wżDu��0b+7�J��㩨y'�ǔ�<�?���Kݧ���='v�8:�5jk�����U���Ϣk��� �b=ߨ0E�@�����?;G��D��H�����G�!��� er�Ja�	��.O�,-|�Ú
�9a?�)�5��T%�ղ		n7�/x�� B�#�ie�s�3��lzyȶ"v�����|\�0a�÷V�Ҿ�w��b��g=g�$K�e�u�?X�)��t�(����x��{�Ƕ������^�S��ҍ�s���>М�z�+��U/
ʁ��@֖��t
��ѯ$���\�'�<m��.�Y��k+@~�t�e	&@�ml^�SAϲJ欿��]ə�6�F���2I��h��v�
���VF�� 3�:@5��S��2����հ���Vy�>Ӊ����,��K)��DPv�ɐ�0>�3l��4�l�{]࿘;u�o�t��m��L�>�i�����$M;!��Ê��c���|Gq�Y�|���y��F�-e��D.��RkK��% ���t٧b��Mskx�k����4(	��-����y�#�EƢi7��/��K�S�Pj��+�N���+�^��&�0י�k��&�VXnl��5��Z\��3���6��/*�XCU�	~5USA#vt��ra�,[oK&k��*g��чP����aT/7��$x���9.�Z�>�m6H�[JӞ@e�+`X��8|����T7IT~]��<�teQ[� 	��������2�r�V���D�����J�����O�5������D�H����r5�� �3r��*�G�~eA�l���
õH�]!��c�Z濉$7�<1Z	�Q�w�G��P�Zz7�d�������ګ�hV��Ũ�\�ee������Rz�2�]6Ǧ!U����h�D�j�%)�3�_�ܳ�����V4*Ȗ`��X(;���Z�l'���Ku������B,�leZ��4ʎ1N��$U�f�����B�¯�{:>�a;��e�:!&���ZU[Vd����p�]�{�W���9��WEM���d*�QcU�/�"W��}B�Sq?�C0d ���p�ؕ�z_��fbC%�����v�ȧy� ��Glj�?�� ��=�BL�U�h������Ynm}hl��kb@�3�y�`�hU��:4J���I\�.��>��E{ɉ��(�����)x���qҿ"�Y. iLt�JE���VVV��|t�)���1F=�W�"��pH[�nl8*�C������=:pX{� /~�6�m�x�sVc�o(�!6�@.M�/#�"�/q�8G�~�R&�+2���{�ϻs���`�I��} �!¥-��J�4���h)n���ĉ�2��{�R,�]�P�H0j$n,"V��?`�do��"1�`mb*�� i�="����ܫT�����	�@q����,�}0T�.���I�e�ɒ�Gzz����y\�!>�C%�e�F��G ���V�����7��n.�]v�YK0��P��w'��h�C�\q���'�С*��j����W	ҍ���Xƙ�����f�D����p3%�I@GVLޮ�g�W�"t�/_�)iPGμ���\@�K6�~�d�ڰxj�ts������񇽳�f�l�^��+�!Su{j	�e��Jm?J�j��@��s)�����1�	�������EO�)��5o���L}o0��/���r!+����,#��t �+�����}�;��ˍB�뻪��ShLz�a4�$됓XO������}��c��{H���f��~�O�9ogn�	"��J1H�^�lc|����wVc��� �j�N,6��P��lHL��@��c����ץ�7�[u&0j9Z�c��5B^y�tWf���pV^���N�_ـZt� �Y,�S��4piq��!�[�>o&<D�(jWe(sKqq��s�u����rk~�4�[/������p�E���isD���b����&+���-��&���Vb����a���6�+����xd�b����c��!�F͢���}�*/�]*Az���k��d����������:t�ŉ����&��H���ʹ���������TP��VA(�Z�xg�J��𶨰c��8����nI2�槟����'��?��λl�V�����c��.c&b`� 9�T5|���:��
-eճ�?'v�Ɵ�d�O��x_��:�� C��St�E�C�*k*�Br�㰂�9l̃���#I�t�5�#Z���(T���"�!xTr��ѷ؟�� �����C*p	�r�{L��f�5� �tZ'X���+����P,����Uj���U,o��`��2V����)���!�ֱ��گ��r������[uE�B���W9,k���n��9��aH�oi����:c�Bw�G��m��:�q��h��@g�qqGv�JGbX(�"-bx��"��7z��~�X��ȴ�Q������~����SI4mǀ���JH���P��<���v�g<A�D�?0	v�ł��' O��0̬�� ��DB���]'�E�5� �nj�(��n���)?M�&���B:�H�{�&ug�iT뉪�ZJb��t�e�rUdB�6�5T��_b�H���1���D��~��������M��_�W�j̻(�,�<�lv]�f�g�g	����AsѢ>U��C6.�B�A���ˇ�B1h(֞�e�E�2���L�=�'N��u�T���u�"0���
Km�]��j��u����]e�QU�����D9T��G E#,&���M�(�yћv"}�/���I���9�+�q"F-�9�a>2�m��C�� T�~��r�GQ����f�"���8(��y���t�;�	~nč��;G<i�P�����[zL�V���3+�<O縏�w�{�F/wB`9�dg�Ȅ�7Y}��y�V�FYk)�Z������q����Q#օ}�� �?������TT�� ���I���].�k�u#�jw���D.�"��_����['��T�����t�@������L���KE�O�J�v��a���7Ob
�
LKc��������f˟EN#���Qz�1KZ�#}���[UZ�&��Tp�� �L(�D�tH�n��RN�Gq�$0~	C	��ԕ4�`������K_��3��-���A�3���GmF܀_�����������E��I(W*v�Y�o�WͰ��*ҡ���x:�+�ô$�2&����a#�t�b�٫�����x���I��fc]Q�E�.�����]_�7{�tX�M����h��N�{�G�%�`d�o�O�	�3lJl�m�W�,��5@Gu?���'������\1<�Z��.q|x=6��ʈ$��V��N�e=�𳩎ݑn�R�6�0X/�q#jQ�ٳ,��R�G��������s8 ��	�5X K���~&|wQB�/��o�@�@�E�_�~������`�-��{{���B��A�Ⱥ��R1 �0��;��,�?��,p*����I���߈�{��%�7u��<G���!;��z��S��d��I�tq>C��d���3E����*���j�ޙ6`��ӭ�� <����O`� �Jh۽�K+���4#���&8��ś>�ʳv�Fv4F%(��?M���sL��d�T�bl �D��/�&�hd'�M�2�0Ft�5k2<G�ÀW{4�q�H[��*DAG*9�a;�OI��<�$e��qP���j��,`������b�E��a<[-x������.t�)[$�r([�?6�̈́3Q5|�R]�f9 í�,������H��l�p�� W��ص��T6q�|lgT��o$O�/�v]c���6".��ϐ���T�"�-���0o5pe�B��OZ^eH�S���9��`X�8DcW�,�ޥ�+���7����g��$���s�1P�y՞�P@;͑�3'�wx��
5��粊.�`� KIѥ]b�4�f�����&�}@?��?����gD,�@z!"",��9��k�7�x`���Xh��ٱ� x�οWS�'��G$[A�(�����ˬ��iMy KWa�Q�g��)=����(=σr�},t�Q#0c�%��؀���c������R0�q��)��S���[�����تLߜ�L��tI�4��?30"��7p�jm�yoJ���ȨVЪ��8�Wxyv��@p�Q���4L�d]�b����G������r�;n=bR������j��mC�D �Vk]j�J��I�E�!� ��D�@���2C��`�G'��Vt�x�/��-tG�XPV�'�������^�����B@�7k��t���@��@^,Q62Il1�s�0㗹@~}�æ���YxL7T�.��{�*���w���I�Q��ۗ$,�b]_s��4v�Q?�� l����(�_��$�v����y����9��8�$1�1�}�.�˥@;A�r�
e
$={�'W��URT���\�Tź�?���Ƒ^ˍ��u%W���kV2���ƨ�����WS'"����X�b�祿�VLq̡�5��	�8��O��G��i�W��x��.T�(�$�Э�2�A�-	�ҞD_��k�j)�(�R��~�"�5����b�B�q�ײJU>���ԓZrV}��ZDm�4��4�rpj���D×$�|h���t�ͳ���ck�CV�3c�UXL]�7�*�R��.��*�qrVh���u��(��R�����wBi�j7�D��1�^g_%�,���kCW���+(�F�R�Z�<?�Л$7{l�>@�Ƥl�����iy�@��ٴrwL�k�^q��$�0b�7�3�l�~8V�w>��l��qS�p�����X�s��9v#�jm=���I�=f��ojϏ�D�����j?c\��� ��*����T�|���UZT�vW�<Mr�	'�UN����A<2��$��O��'Ub�������;�
h}sU�a��a����_���J�c�֑���[�'��$��oM��w�&�O_"� j��o��A�T1���Y�`�J�z�<c&Tq�9E�\2Ï�����CB�ˬ��$@­5��T٦��Z	�>����\�k������o���<,f/r�˅�(�<͆v�6j&�-5m���:����ǚb����W�P��������� 9�MsD�#xSg�oϴ���=����T��\���lG|�b�d��o�m��_<�7����#�]t�0��NS���{��	�{�4���o��irБܶ@͘Z�������ve.+��7�@��d�ε2J����h�{�'�ħH�iRGUG>`�ݲ��雇�tӝ8ƈ��oM�8-��������ه��x�sƅ�,\������5�.�U��)��U��>�'���nH�Q�m�}��V��ɏ��L8B����tVF(BQ���0�20��GUR��uֲQ��dhBN
�"���4���bP+��H�m���4m��B�e��SŜ�����59�Al dI4�m�RH��jѕ\��Q;ٞIAvb��X�5�q�-(,N�|N_����X���Lk�<(ׄ����p5�3Q8yn�g`O�9�Vݢ ?�i4^q���MRE8*
C;m�A鶣�3���XA�o������qe �z���A��^��#?v;�%*���+��xq�Wd>-\q"L�,�Ӽ�C[�؋��6g?��Cy�6޻X�7*��v��]{�T�����vh�;݇��TM谔\�����PQR߽q�ڠ�܊U�k����|��dVJ��o�	Ӏ��v�72��2'<%�9����3\`��HC=�m�瞧�уIN'�fT-C��N!`P��;�9	��'QE<޵�+~�S��`�V�4����M�u]Cg��"L�~銟L�}�qkP�<��StIMO��<���6c���n^|�wV:������ڗ���T8���p��Q�h4F&N�kL�m��uVJ-v�����4�ֲ��6�sX��O\���5I��2 ���������;˭4���7P���@�x�)`c^`8�>�ѝ\!D5r��\.'�#�\m��X�;�������1�R%�*�{��T&<�t�a�Y0�H���z�9ڹi��M�d�`�M�%�qa��f*�E	G~+�Jʼ	aʏ�>.r.T��RU�n��i'�3���bJP�Wǰ?h��QiRFCG��"�I),�K�K��7I����p�R���Nb�Ӳ�;��D�5/���I-.����0��[�2y(���-��Z@�`�#GuTjK<���v��b5�֌�XC���Y����h̤���c�g�,�XN��B��������ЙN��O�:�1���]�#��h�;|7C�,�R�7�2������B��W�xQ�4�_�ZC+�(Z����H�	����6F8�宇,Ƃ|�n���p �X�P.ow��g�vQ8�7�<���l	o��8�n�k��<���J&�8rZR�0����х��AfZ~E��4 �Pm���zCqn����ʋ8�}^Ã��QJ���K�b��Kq��X~��:j��sD�
��Ź�5#0Z��m�
d�rUُ���=w��,��ȝ��뙱��G�?��ݝo��R]�u�n;��ۅjsq���	��0�̳�������{��
_�p�����%-�*�s�b���������\<[ ��Yț0C?ϫ?���X���m-�e9t*�\��,ƞ�����z�7�{��r��a����/dW�E��p�=�*��MW���R�T�}��O� )�%��Ǌ���@NKwc�rv�!������V���Wg�u��^��j�Z;�93�f�z����bRD�[���:�.��ڄ'w����ü�E}X_x�R�QWU��� Lރ��]�Og�A�ƑcTG���2�U��|XIx����|P-*���m����B��T�����0V]:�IP:����Q���9��:vS2����/h��>�r����^��-���#vm��n�`6�)�W``�;�N�a�C�@zrF�V���]���O��6Q&R�*"��9W�?8� F���|��z@���H�%R��ә�:ߴÏ��Ŧ4K&�`(yY�H;b��Ni��|	�b���3��IKPn��EWw7�S�J �L�_$N$�����ؙ��0����_|x>�UY�4��K�>�U�\=3=��(W�T+�OC��V��r�2�4���-�T4S,�Q	ك:ئ*��4��c�De��wL�a;��WQsf ��x�W�9�����^_Eu�s��בl��L���Z�ů��q��r~��7��B���띷.��� d��5q.�b�/��%ԙ�-��8�\t��5v�$���"]��"9��i�J��w5�/�"K�`�[N41*�2��G�����5��{�L��B�?��?^����C~�_CKÑ�4��}�>��919���>��"|�B
�5o"p���"Z��Yh�1�>}[N��Bvp4#�`ľ���E��oy��@�NO�ǐ�Sg�z���uf'� x"/��[�=��<�"��(�|������Z��w�MK�u���:t�;�I�s�����F�8嫮@�滔��2���2��s?AZ�8~���g��CkH(`æ�X:~�t)����l/g��#�>�,���O����E�����:��M2s��<�F̕������&�w	ق��f��̤*��M(3Y�s��/��j�C�3��Z`溜����ss��?�oAwgRt�R�}!qdi�x��aP�1��
�d���O�w��ӎc2r u�D���~fx>��b@uy��
j�Lv����Q��<%(�����	�3y}זΏZc�X�7D"�t��ʮg_�}�{�+��*�!`���^$T�LHE�����K8��?��L�	�rXG� 5��9��m���،�\ќ]��z�y���\�"&]�
�ԍ}a�O����/�}��}���-�ۚ�ҩ�7�{����H���Ǿ.�ә�U���V�Ϛ݄��I����X�>�YZ���Q�WNWb�DА��׻q�����^��(��rz�����C�,��}#5��W	4e�����1肬;[���k�,��F�y��m鉕��Ӵ���80nް#�Y�,�x5^�J���&��2�v����YY(�P��a�<Nv*�`�G���=C��� ul���������0��;��/m�����<%��eR*�)b.���}3���ܷ,�Y;��r@��|KҦ�`���!�wn_���!T��8>�R��9|��"{�I:t%��ݔ�+����8��IR�6	'��B��N���d�+F��1[��z]�s�̆�?�W�b<\�hX�Z�����d�XWr|X��i�H��cd������%N�(��,b�Qy6K�}~�2�޶ߌ�$A�z��7�ξ��|%�����c���"��=��]�����Q�ѧ�v�8����&Ä�Pt;��g3I"~��N�b[���G0�2{#@�1]�.R�%�D��V�	[SN�{x��%%w"!'�¿�׈���E������A$g��Q3�����I�1��(GAʁ�P��c�%�_y/;��'UW$g��ןyH7G.#p��!��j}ps���܌���2�#�_���P��{Z-��)c�(2~�14?1�j�(�l�~�C�'+�Q�y��R�57P�����T����Yp=��U���%��z!��R�RD@����b���>/��4�Hѝ���{#�h�H~ET���ؚ:�#�@� �-���)�mDq���F�_���N!}�a�O?�g^�.�R�����&fj	h$����=�y���W��������F֚'	*Q1�������8�hg�E���qxŮ��l�m+3�R,���"�>��̷�Io�Dͯ�T���Y+�&�+O��uV#q�>,�ھ7�����K��U������˂D������RЮ��6��R�vH�%���S��q���JRAT�N����/��:OvI�ȵW�#Zz�`�lz��<<���F�q��Z�S���讎���|��ϑC��:67��Wy⤊�6��b���#g1KQ��jWI������v�F���b��Iȑ�e'�j�5C���D���	����k���@��st���OSK���
֤΄�.,�&W��>��Z����I�b�u����mg�f
5�~���f:�~=[~�z>��Ja}�A��ݥ0�Dl�l�� o�F�W�+lU�F�L'��d-��z�P�!&|��o�����3g���u���H��B��ol����M�'�ԓ�60]�}�-��Bq�W��3�[w���2�$� M\]ZL	�*t���!�;غ���Q@)r�*�0^5$�ç�I	���؉8&V��l�qs���X�_�gF�n/Y�Q�XЋc]�6>t�b�B��v_�r?
��\��+
�
���M%H �ֶ&��!+�wQF��x�=���9��`F��T~�|>��Ā��(ȿj
��ԙ*�8��<�:1�C'��@ل�H��y<)3 �pI�A:�&���ӢCOLAp��|���(�v�|.\Do���4��eU���5@��m�� Bf���/��T��&��+�j�3�@x��gH�D���u�E4Pp鞍pyՖ�G�����c��+�|���]WnG����|��.�l) �е�[���|#*9�Q��?�QE>��Z��+�*I�eqo�*�
'�r�^rĝv�~��xe-6�~�@N�x��ʐ?�������37��T;�b9��sM�������=)�{y	��$����Y�{&5*B7T��^�:U_�)���7��m=�d�ԭ�3-~��ì�i���cp���
���<6-�����k^�,>����R\"_dr��|���I'�e!�O���\��ߥ ����������$�,�� �0ƭ���pd8����KCQ�vrt�|  *��%��F�"=
��A��[T�xNٕ���,�����[`��xv�kQ� ������v�	fSj�Ŀ@yx��q:y{�ߕn�S̍v��(�⑍V	��M�)���'�7: ��j����f��F�(��{$�ɨ]�[(�-zy��WmK�����?������:6 ieZ[��z�V>X?;�2����R��W1������)�e�#������7��Σ�n����
�'�EZ8�U��S�q��J蓃�H�9�T�@�#Q���<%�f Haz&�Λp^�@�:�C�5GE���on�����x��Ǯ~�݀�;��?���b�5)��ٵf����1BҦ���MW�\�<��W#���N%W��*�����X-��_HѩX��]ɐ�"�K;CI�T�9�h}s�H�I�rs&��� G\�L�0�~s:��dQ�f�a�r��������M��~�r��϶Np��n�;�fR\�� �	Pܼ���T��$oZx�'����c1ֺmF,�p�;8�:�sX��V	2���2xz���rS������%���hQ��h�*[�	sV -A4	��R,�1b���pF��ۧ�	�=��JX)��Q�r���bGx>"�8o{���%#W�ÒT��ڗ{8V���>a����ɐTb���T�� �'�R���W�^�IE�G�#��d>��x�]�|&����`<{�2I:;�̎ za���/'z= �
���RM�мY|Eǆ䎪����G�%����0��)��r����mGJ���h��#�?�J?֣­r��T��)����'��e�.��."[��`��p]�<3>�K�Ւp]�o��gc���F��&\�Р�����;6B�@��׍:PRfo5�3<vv��-o!椰*\	[^��w��%��R���H;�0�_/��)|�F�
ڌ�7H*i3ƪ�PX��>�L3 �ꛔ�vŇs���@IJ=��,"qH��qS0�/L:8o��#��8��	�|�R�x6'4�]� Y�%�s?�������}4��jc�|Q����].4������f�Z�b�x�ZE&��	G���h������M�D�N����h����Îa����L��~yN����|��g�$Z��.m��L0����ԴJðr��p%r�dA\�&i�������-���6`�Ď��t�.A�ⳙE����č5�/%��8\G��\\.���)�П])�(nl���
�m�f-�a��(�5�A�6dri_�] �'s�]Pқ(4��.��\_�-�v^����U�PNH�_�$�/W�Q�oW/��;�}~,Q��*8�x6Pf]�Zk�Q��6�X��YA�b(�J�O*Y�{�dTf��5N���B�����܄; 6/�綱ǜ#��(��6��c�X_BCq0#�y�]����6#�Vh՗��o���}vIc4mbO�E��*�L��?��& �o�H�k�35����C/��Y�GMv��x��"��hoi	���B�0p,�wf8��C݅�;�y�>�\}��&AP���_X�7���;ac�b����?���,Ҁ[���ֺo��IN6�}�'���>��b"�ӆZ����C������ q��pL�L��i�8�7{v)���Q 7|Ə;��J�E�#Z�g�Qt���^��N؎��8�q�K?m�R�!`P?�7��obĄyAY9@]�;�M'NP�d*��:�@ �v���XI�����]�ίy*z���Ϧ�1����o�DL�yk�܈���薋ׯ�_���\	I{�����hi7��cH�#�7��Z��J�m�:Ɛ0�+�1��HT�	�eGkE�N�����Nŝg���<0�i�X�,C�����P�;�Ai�� �@�?�ʚc�օ/vc�n�3�-�F�(w��M�>���sآ+�w�׻����:�R
K>��@\��+��\�c�<Ϭb��$nY8��Ӵt�,��%8�M!ڳ6;�"��$�n��X];�5���v�5[�z���;?gQ��>ϥ�Ϣ�1�v�h}�d[Fn��:O�\-�U������i�0�*��W��;4i}��D��$8jt�+G�]Yo\b���Hz�Om����/�;	.>p�?g���n����3
�X��V�țA�u?��e��|q�Inʬ���dbhţi&Hؿ��on��T	���?G9�{�Ā�s�����Np<S�F�ژ�.��������X\���p����iR���
6��Y_�m��/!M1�ǰ�?�)�g�)��<�1î�
��s���wn������(aU�4	Г!��S^��b9iѝ�{j�3��	~�/=��w�l�$��X��Z�~'Ca�5;�e�0	����a�n��ؑ�ꉕ3(z@'����^y��zYɒ��2�H+D{���7׭6��m^S��R����H���81�1���{�$���H��O��}�D���6�Y`�h}#��g����׷pD�� �*�oJ�Γ�+�(T;V�ç�o����;K�	��AڻW�c�{�ũ���P/O� �;���k̾BFy�V�/ˑ� �b9��C�d%/fL-gp�m�&�E'�!ci����;�jT)xaZ-�9ZA�%9���a���6O���H�ϛM��i2��Vr�DuuL�SԵ\С=���j|HHȻs���K�=��� 3���or��P�\�&�ݱp���q7KѯF�۵�'|�hid�<�����6�)�;[�-G�w<�K���<0]0Q�O��U��^i+Bw���1�"r d���!�w�.Vg���#���׋���r�f`���;���P�$b�w������!By�\��`l���(P2,$:K�NR�,�UuC���'��ѪM�$��,�o�_��9��Qa�8��}�@�;���J'M�_�d��3�ݜ����(<����.�?4���C�Y��/*R��32m�^�~�K�T�0m�b@��D�#07�,��`��jD�D���Q�rǍJ�&)�5�`1vU�Hߙ3,�1������2OQ�;���)R��X�9����G�eM��ޘfan��k�������V�/w�0?>���ﶷ��`v<��3X���K;�HX�����7Y�N��goV�����]?�(�R��v%BO^��&��4�I�PZ���T��h��?��.�A�g=��M�p��p
`��)jA�r6�P[O�$���1�m�6��(Z��7���o<�w��"!9�����>P3���n&����J� P��"ݡ� �OW�Ά���׋8C`ۗ���[��T�?n������|[�����.��އؽ�λ�\��!|L�k���?�{�+� ��V���*�T��ʇ�C|��86��2e��֑)U���-ξ��-E^��Z�Gwg[�k����D
;/E�F3�sQB}��A��� �.A�����>E^>��f+QG�����~�t7o���T�T6�"K�>�*��=9����@����j�Mz
�B7`he��h��zd��!P�[4�9\l��d	Wx*|���/a"rc�Yf����>�@t�}�0ŝ��m9�h�	�G�q�1��p!i�-�G��������_O!�e���� �%�á1��3���47;k-�u"�[�_��~��,�p�X�8����c"�:�S�dt�,;=��<��X���wy/�C��D+.�񀯹k�Z��g�y�m����J����|�ȩl��˭|Y�N��k�Ţe��J$��/����c����>[���^�:��*�c����Gg�f��q���vh�@v�B��xX܆,~Ѻ��A�)�i~� }��L��o�ǐ_%*��OH����� �8�x"'H���7��g���˽G�\�:�v�hq��T�۷��=�al@?V�]O���5��	�4�#�@�A�d�B�d�!���]���)u�LPl^EW��|k𾍀�$�r^!�6&u-5����N�I g��<;�0�S���h-.W�x�&�X���C	�=�U[����SP�!�������Y��0|�X�m��Ԣx����7����!�i�{s;?�������ϫw?�!�Ww�iP�2N���}���Z^j��s ��|B��I���	ֈ��n%� CD���E�|��)]�i)����ZB����Y�H��=�j���-�_HGJ��5c��e�C�e%���Ƈಫ��B�@^���U�]������{Q�`M�w@g�}�͒Tqt%��d�v|���ͩ�w	���r�e8� L!��B
E����H��h�P��]O�Y�'���O���]�1��"E���2�ݰ�|�![;'��5�lƤ^��e���F�S��r���4���D�0�~4�����E��<vS��k~�AFy�½1�̍,�=���:�A�yy#�1|����	�R@�T�0&GT��4̟��$?���+d�F^	�9�y'�b� ��|	���WKڛꮕ���e�{u�\}Gl�[*�6��O���"{�5M�A��YUl���J#�d�g��w
WF-K��F�\C9�.(G	<�oc?
��м�YL"J"6r�pb�R9t�Z}�{�u:��B.G~�i}���$��z-+48�$�h��L�<.��9�g,��?�,�Ml�L��U�8�,D�O2�,-^I��'#e�	^x-p�C=%�N_Բ�5Ї�Ү!��((1ߡr�����7ոY�o�ł,�Uk���$�)+#%��}ӟ�)?V%s����C�j��$�[�͍�:�g�-�H-���p�����nݫ)6|C�q�- �|V���'p�D'=2�-�M���Yi+��i�n�E�q?G�uLTZ��~O�ْkje77;�#��b��wUIG�s���DZ�evؼ(ؿ��h�D��/; �]�Ն�eZ� �*u�A��wڰ������a�?X�σ��N�ɤ�s�4@6�*�5ʄ�y~��g��!_gq��a�(��bە \�H}����Kl*�WQ��#Jo����<�{��?��%Ry�y�Y�%�_y�ע�%�CQ��Shf5$u�s>�
���&�'M�U,#Qm!;ڦD�&7I�/��eqs�?k�m�$y�GN �%G��-7ff>���xv1�r�mg�_�b��0%�R���g6����V�[06�↗"05c] �Tp<5�:כ�;F
��O3[���D���@tjb3ӓ�GQ��R����e5uWV b�A���ØkZ��7Zz���H��iAR(�� İ#�<Wy"�����r�� �f�m����(�q$;/�96�忻%�D:�|�<�	����>��D�`I����-@��:��ϰٱL{&�bL�q5~#+Ӵ��t��A�~��h��@�E�z>��V�V��*�*�}g|�����xf�B��o�?����P�-��G�������8X�ʡ�w��ϻ0�m�5����t��;y�kk���5�����ɧ@4�R�j����m� ��Z͟W�*ңΩ�A&/��[ ��#�}F���&3�@��!��'Ӆ!�1����t:\;�E�}��oy$hM��M��4�`�HH%��HR;<H��T�Z�)a44���|�O1���Wպ'��W�t��\Q�Z@�#׈�'�D�E�L��h=����WZi��~���1�T�n��t�����<��P����h�
߼�����Y����܀(mb�~��Y/��>l��ҶL�SSR��.���;K��?�S�Hq^h8?1؎���y�g:����1��'I�U�Z1-�o���Ĳ�� ���G�	+��gu01X� ^�|Q����(R5��@|�fkH�K[�OB��,ja��B�ѬF;8.��@6 y=9����ZR4�'��#K��D�4l��~�u������l��E��k�L�fs�8_*���\�L���ޓ3>J�[�J�b!$+���WO=���ɰ����e
�
�:Q���{�V.B!��"k&Y��D�����L�_q<����	�&L}J1gjJ���H�b�+6�$_@gp�ng���GF����pZ�?#=]�ƳE�%����ƕ�@¦4#�:��1N��ü'nDM��Q�0A��5*���,͡	����/
~:�A9
G����;]�NJi8�4Z_�/�X�F��������������%d�x5�\:�]�Q�%q��VC�P�u,l�u� Lz��$��;𝾻.A��x9:&����[�yf�
,�qX�Srx%;���������2J�T`�����=+rG�ѧa�ڶ�g��E�����aL���"�l�m�
���<�6&i���$mS���q����6�j����G���0�A�p��N��yW
��V��T��^�`��R]����?nɓ�ͮQ�VTF�,vaP tZ6)���{s����\{e|���K(w��[��-Z:Vl�G���5sK��p��Dl��[�E�WҔ�ӆ�
�@y�����.Trw�ȿ�O�$-�n���h�|B�`SĆ���E8�Ŵ�1/��܀Z��\ioQ�L����=Bɹ_ox4��ξ6��>�5�L�@���̜XI}�a�:	X��
��m�WN�ecB�3M�g;$j:��j-!.p4!{,A*�WښUχ���1�S#�r��2b���ND]oa��v�"	���{��"�{��49J筞щ&@��ڰ�׺��.��n��<������W=�2B�TX�y@���U0V:��yiw�-դ�~�z�7C�����\}PO�j�)��z��s�&�~<�<��ZG����{9"�MVxSA������:hr�A��-R���wр&Sa�Hr5��;,�Ϡ)���i	�6��� fN��	�ݾ�v��MVBv����4���5�W)hQ�n���a���(K0s�������24C&�֭)��M=�jD� �MV��� �)�k_�]���e����!�����n�A��� �xs�
xH!Gcf��IQ�C	t�qd����n=S������:1�*�����m�J��J|	�F�D�T����̡�����m	�Z��Z�uK���	���k�}?�^�+j�B�خ�
.��ԉH�������r
7�?P�!|�T)Ĵ�)��v8�|�r�f��QXhp���J(-�[����7�Th��uC��Q �g����arR�	�XLs�r�G+�l�᠑X"
[m����u�Pu{�W�ǻ�Z`�\�������is�OQ�|_���;rc}J�^�{�Ǝ)�oW-�#�]g����K8q����S�T��թ��RQJ���8iF����n��|	u�r��a
�V��-��΂�� a� ��[�ōꄇ3�	�P~����K������dr�^���K�ݦ�z�v��,�fO����0�U��+�ld~/���LA4��̨���G�­S���v;sڲhfj����C0��b�,Nrw��#�2�cKÆ]GT�Z��07�y\?m��K�a��YeK����	<��p�b�
��^0b��[F�� dJ�iq����UY\��Ҷ%���;9���/��~�
OEH�%U.��JZ���Wv^V��{�w���3�{�GP�Q[��Hs��W3����ނ���s��3+��4H��f�c��9D%��!�����;���K\x+����$k6��Ơ��ySK��mo|�p�;2rʙ�yq	%p����;h���X���V�o�,^}���������O�l�~^u��~Zi���6�Š��3ul@-^��M�H��8ƚ#%�-��t�\1� �}�'��TW��1�΁�,jb�vnj�v}ʤ��9�?���a�P��/p[��N��8�\]6����L��2�mЪI�}�`��S�Q2mS��j���)�ˏ�'���7XlUƱK��G�$�HY�����VlQ��j��}�"���eY���n��\�g�|��x��
�E�w�,�QX��F�;�1j���_������l���n�| -��'v�y������n ���&�ha�KѤ����O��Yt;�C���@ɍ��!Ѣ7?���M&Ĝ���$�#�2Y$y���`�Z��i���c����v�yFvCM	 [����u���)���M@JHI�ި�,c� c����ؒ[��m�D�h�Ԇ��5F��'̉���������������Q5ܮ�:o�:E*����Ep�F�k,߼�Gr���E䗏�=0�'PO*П�D�7�3z�����<�ߪ+m�/�S`.��^.�������]y|�!K5L��(c��b���}��?��4�j%4�c�WLˀ��� {k��ھ)�9��0N:X��,5}�͵�������A	W{��W�=��q��|��}�ڃ,a��a.�ھ���B�u;�$O�֏�֫=g��$�h����
y�6yY������s?���	�c���jpQ����g-�H�����g�7��X{�y]S�������wKL���x�lm{���!��ݩ	&R��[ѣ�]��"�.#�h�6QT��<���4��v�։��BB���7KZ��|���t��HCm��ʳd��ú���l�� ��VR�V�E��&�o�=d��f�5��jy����"���q�U��|j��v�΍���I;�f7��Cϱ��6po��<��Օ�b#�.�*u�.�}r`�c"���x'Pv�?�8���P�Y�L@
)cd��� �v���hoj��ٲ򂺾iן1���=O�ݦB����x66��sp���M�&cȰ?Xl�j9㶾��xv�=��a��S��)h������0�y/�M���#wJ?���G�cLC$�J����� <�cJ�,�����wXm`���E��T�vvbwjp9�i�)G
k��y�g�w)����k�~���%��F}�.�9TZBߥP��x2c��w��~;�wʢa�8t � �č�^� ���z}��i�A�������;Q���Ȫ��h���l��B9[y ��z��<��",J����q���<���Bn4�B̢�����a����&m�v��鐀�0��{/9��<E�f��4�0���b�O%��d��9�J��ޡxr�z�/�����6'���8�K����@��!Bv?n�8Ck��9��J@X��(�2#�e�X@	*��(����O^�I�"�W* {�jG�)�gh'��0�����Te��"VP�\�|��	���A�7������?�g��S���5��$,$��W���߭^g�f8U쏸�a��V�B4�97d���Bwgh��E�|r�KS�O��'/V+	`|�+`�YJ�����f=@�"^�'-�p�'m��zٓ&�<��
�	ߖ���n���^�H�d�����[� yС%���>�d�l����� ��D퉙(�
���={��b���e"Qs���ˁ�B[j Zŉ~�������E|�]=?��-�s, �#�\A�d���;r�[�M�$�!	a�Z�(�/�l��
i\.W�䥒d���HGK�0+!ka��D�'�V#�vOf�\���,�,F�s{κK���W�[�1���$c��scy�ߋ_�>]��V�.7Ƀ	�6�U}f�!�����:�&�a���a����.�)�]�I�H����{�;Z��z`mU#̪�n�������K��݇]�p�����Et�5N��F����ܥ�@U�_.;�<4.k��G�61�>@��A���-�Yd�����'�n�և�<3һ�������������{:����e�Zچy��5�8�Ul������l��'&B�Q~��P��NH�M�]:���fX����~���g;�9/�N5w��y�����	 %s�J.��JL���2�<����Q����քD ��.7�k��;��~���vB#_���4U��Zc���+6��޹
{�f�����A��,;��?8)9�X�ކ�v@��inđ�v@eH,,��iJ��gp/A��ظ6	c�h��T)�vZe}��:c�2r�GX�:Lɰ�L���I�ڌ�$�V��(���x>���H��S�cg���������)'�ZT�	���5���]���ݲo*XD��?�j��
�}sΒ�J�Z��@��X 7)�4/���b�D�3�vc]Z�?d3Ñ�P��l�8 nB`�b��7��J�����>�z����?&]��>����3��d�A�^�H8µ\ �R9=����l0��[_g�m�<�C%d��e�x��4JEa���eܹ]��%Q<�Jb�2�@��j��<�o���@ ���!_�Y�SN���k؊�-
IAc^���E�g�^&�v��x���yf�*L�Y|MH��J�k��	3 (��������h��<;f�~~�2/:�k��\�1�&�w�BY�uU�81+d�����ï�SteC;�Ѽ�0�`v�OD�-�ԁ`��d
�~�Q��bA��%��f��W<�WN��j
���`"��]��3��8�������A�A������ �@}j8���@r4���?{�Ӽ(�;���q	o�qi"��������B�F2f�qk�!x�:0�>�?%��hVEC��Wb�[w��E�0����
Zt��{j)o!b�R`5�u�e'��i/��fO	wA^�[@���\'(��F�?�u �P 5�2K1-�s�x,]TV&�L0�%��%��fJ�wΡ���;�N�h�ޒ�P�w�Ӥ����υ=��k��8����T*�i"�+[�q$v!`V~�Z0뷏�'�T��k�5�R��(�m�o�F���tz�����Y��g�*#Vpё�H�Ii��������|cg �,N�<X��*�e��03����m�ہRB��?R3�|�8��;����@Кf����C��_-�[}�Ѡ؊ۜ���������{��o �`��0�:��g2��o7�FP�5M�B�E��� ��8�&W�>7�Y��+�Ih����lig���L�w�5�ul�� �x�Y~�d׺��`���y��%
g	H���z&!_+���/��;��]I�P"����	j�e(su�7i�01���+�o���(�Ժ�7���
4���)�|��U(ߟ?"lQx���ꈶ�Z<h(,]~��ͽ4!b�\��t��^;U��J�؂w�Е�6CJ�-@��g����u˚���S.�
��C���u;��K:T]�Ϡ叐�AS�o��"f�����h�h��0+��3��3��;��l�)@�<ˢ��)�8���S{����D%iյk���m�G� ْK�]�ڦ=�Ҝ�y��g!f� �;^r����R����l�K崬PH|�Ҝ���d*���i��"������]ߒ�g\�W=�1��Y2��@KT��^j�h�!ڎ�4K��x�M�']ZeĄWu@�a������>�ȍٗ��'l���b��g��K�c�i�2"�^z�|u�� �9V� *ļGX���(w�*v�-��U&�P�o8��{��ԓ�I��.�E^f�pY��%;ۚe�νO��%�\���<�׺f�pP߂�����W��!Ä�(v0.���⛊���2��0��;=����'ew'!EM�T`EH�0�2�A}3�T�����J��6�h놨�x�Ó���0� lR���z���O�ˍkA�٣8��<y�L/G�,A�[48a�y$si��R�������K���ɿ�٧��^O ]�D%�w'�:X�%Z�n/҇����-�Qv\�>�d��B�f<\�`�Gr�vSpq�t��]�ez���t���"2V���O�ܠ�x�~�xn����ni���(��N�w���Lw��~�6��si�i^K�ο3eW�40�.�'@ׄ���'Ju��:�A�Ctzj�6��V���z�lW%.�������_�<`�OmPM�7/�� r�$�Q�a������� ��aB:>*�3!����LB�SQ��X,���Zl?�ۗ�0�ې�
�}��p�n0��Zg�t��`��0)� �O�qo��	�������|P�@���6}{~Dܺ����	�D/�7�6�艞}%�똡D��lR����6��	�bp-0Ҝ��B5���N�k���ї�<�a��u9�f�����禝��q+A���S�[F۩Lr;%�Tf�~)+��={6"���7��b!���.�Ǩ�-!��
���]������ R�������N�#�/!	�χ�jc7Sm7XL��<�t?�b��;�%�H���ef�@�2�B.IK�؝�L�(�D��ˎ�n�A��髦/Q�۶h�I����\�o�/���wC7�,wW�*���}��ϡ��C"�6vv:_�O�b]�#z�.2��.�|���-�Q�ґo��DJ� aMU�J��4���~؜'��GI��&D}˿�O���4�})�Th?'��rF��@}-VO��� �@���P�Nf�,��6�-�t�(�����z>+?b;8Hho�*��=g̚gܠBnM��؇�����P�i$7Ӧ��Ъif;6?�0I�!��KZ���F�bH����ygUu�LT�����A-�Q�<�Y;����IB�:�_: ��HYY��/�ҿ�3���ghkm[�u&q:X�$yfM��X���Q�y)�Q���@e�uΰD��Z��w��`?`m:3J�-9�JYd��E��kD�gϓ�'d�L��EC̬}��k�g���x���R��#ޚSv9�s�v����.��q֭�=r� ����	��� dZK�i�+U{hG���Ҥ��'*�4�1�����G?J�̷���ȳ�Ax.N_���d_���)r����6�|^v�jb����7B���M���Af��?|@�Ap(6���N.���xλd@��������E��5����mZ�u�k�&r9�?e1���}	N^��U�����NѴ��.����H�T�?����R��iּ�s�.H��S�}�l���u_}���%qX^�����E��]y�g�.�*�k�ZTF������a�k�\���惄��Q�qU�S�mBj�B�z��q�_����9��-:Z�8N>i�����Z8Sİ����P��߶E@����fu�Y��;��VaM�z\u�##7�Q�x��FR.����dF�ۣC�h_��a��0S�^��'U�8c�r*�#�7�I]T7�R������ݺ.��J�xP=kr������K%�Ye�����<���D�A��ާ��	�xU�+�-ܗ�g�}��˳��ɢ�R���ɏVx��L����'9ms��)��FM������\�V|�����6tɘ���0��0i1�@hJ�Q&�Y�i�	u��q՞����ɬ)!�J��j�|SUaz�ñ1'-���w�q>�1n�%�<��/�5]�M[l��3��[��(z�!O4]
�y]ZkU�rʦ^��C4����/���2/��]������/j*C'{�Rv�H�Pp�s�[����//�,Ș }Ei��uY��<��.WP�1� ?��7Wz�>�ox�%<����������#��1����e=�j�u2���$��ĥngi͇�������#��q��j���`B�9�W�T>�]��S��_���� 7�@����t��L/�Yn�P�F���b�e�ZZ>�@=!�Q�ً�q��WI>���P�ߦ{��@Fͥ�&b����!��狏�H���<i���d�����Qܴq�k��*<�)�t�1��]��nTv���3�����Ɋ���=?f��{p�-����(�������u~�igq&��w��'��'���U3���JA�;k�GM{������;Zi�;<N��Z�3��-`�]j�[!5����u{7���Hx�9��h��H�}����t�wp���ڒ��z�ؐ�z�O+4B�,��<^��혐���Q�LW}xV䖐��o;[D��\D�)H�C.����7^�=![�)�������!C�X���-@"�����:���br�C��@�F�°wQ]x)�
��h֬
�!�؟�Kj7�8��Q�+ߙ���wvW��Rv-,K����=xM�%�bґ��B�b��e�!x�3��W�m���r:�	ĭ毇�B�-Yc.��y��ܥ|�4�$�����B���TA9�����`FplT�@�vjV��zC�H����t�ň>��
w�/��j�7��lK3\4?�hZ���G_�H�H�n��,���0��	^R�b��>(�x�ް��]oR򐑘m�<�A�+[�d�<c�E>e�5����NN����ȟ����2����wS"�0f���n�\K�Ē�x�.�t�F�
n�����&�E��¡扴 y������n���RD�E��͙�G!��I�V�;�mw��^����Y��S!˾% (��Rv2t�����
M9��7.�~,�`A�*�PL��D���m1�O$H2=�r��D>Q��H�8�,����Wi��R��!�J��g1��90�ɨ��:5��`���@�̐�̚�5ʀAAM�=mF����KF�5u��%�(l+}���\�-bT���ѕ"G�T�[a$�)"~�f�?(�)pj��gP����s�>�}?ƔX���k��bGb���Nn�EG5������!4 ������{=Ҷ��_������3�2<�j]X���"�v(�*�)gXx�m�"�����~/�ѫ����m�`g�}3����G�(���?PB�3�ŉ��J��t��r:�SI���)�U£ �`��5ѿ	�g�1q��'�i��x��\,h�T�s����[�L�ܙ�5��k����]�N��38a�|��UR��u�������~-(-T�<�M��RTL�������i�ڧ��s!g{��u��Bz�l�0���-��m��]��h�<@�It#��7h37����윙��,Ҹ	DY?<��3�-ug�̣mY1zw6�V!S>e..���|^@<Z[=D�� >��Vy���k�^��/ę�g\7�g^4/�6Y�˻#	�w>dZ\rLg���� n��Z�8�"�N�"aA!��G�&(�V���<Th�ݫ.�`�ME���eξ��9�M2@���nJ��BA(��̃*036}c;X�IQb<9�.n��8�	͑p;��Ү_�e�=��X��C˔��@t]�ꈕ�i�"��0F��r#��T��x���10��5p?i_��K/�7b��Bۣ`nHX��<r̴E�\D��RC�ZBR����R�6*�rV<�4��?f�2�^�I�d!�^�ߛU�Z_ğ�SoT�׬*��÷O�t����T�*�U�)FDN �n������C	m(:@�iơ9�a�~P����,|82�e�N�����N�J ~j����-bP�A��-ƨW��{���pH�tb�$D���K�c��|�����`A�Y����~��{oM�ۄ_���A«��h����m��&�߰L�����0L�8o�����,���
�B}���zǁ��%�ɯ��_ٽs�^W���v����\+:Fb�A���]����]��@�N�@�� \i�+w��q(��~���
ێo�@~�.9����v��_*0:W�K{��{ֿ,����Q����Ϯni����ؕJ"O0g14�ɞi�N�&,�[��፣���E�����pI�G7Ş�{�
�l��%˖Qi4��&�Yx���N�F�������F���m�|��Vw���|����J��*d�r[@�;��R�I��&���x�σ����+LxAW���IPK��<�/����&��HlcwNv85�c��i</��ӢY	V��!���]zmŮ�UӲǹj�c\
@d��o�������r�F�L��~��l;�M�Mg����
L�cѮ: ��bE�{�7�����Dʧꚓ"��L�ީt�4%��5��1���|�Ti�I�ѥ�'dr���p����Ґ�J"�V5� ���������6�o���ϵ��R�>����F~�ABM���T1��Y|G�q{A��c��/g�y������=v@���jO�`�xjN�s[��)Wz^/KE�U��[#!�4l��������$��7�gU^ўD�ݹD���cf�k��dх�nKtˢn-�.N�dU����
Zer���M����q�s�TB�YG���Q�@oC7��>�=��~����j�k[8��B������H37kA�:!�㘿��/����v��j��ț{A}"�<���s!@:�FE���*
����Y]Y�h,�ŵ�n���`M-��E"�*(yӓ���9Jy���emE�>��d�A��%��4�����ޚ����QK�Qæ�&��*+���T
K�o͕���o�������e+rb�O0
�YcVŨ���e�(R�44N䶱���=Ծ��f1P삡nF��iu�^����Wu�%�ʢ�lFJ>��`��Q��'J����h����/v��D����f��_�+<��w]Z�z��Zu���<A�]~d���8�7r6�0̴Q�Hd��?��O�<��r�_�[���V����V��#S��������t�ь0~knc�
�+��n��D�ć�u��=���p5la�nl�!��3�hh���`��r{o���:��q`���}����k)��w`*&�F�+�Ơ���t0]����^ti��4���7�g�WJx����vF����|�X���|"�An�ofw��\�&
�Qb��/��o`�GuE�5A���%�	<O�0h�k��]��M)��P��_�/������!4��-b���!�PCZ'���g�>��B��g�������^�C����sZ�7)��%�����F(4Z'�c����L���R��5�2@?�j-�Dᶮ���L~�.��b�X������wx�^p���f��j�+��������O�]��iq-q��_~؄�E<���z�>Zd��$r�IY߆L��ST���Lbkі8����#�E�����@�*B��3%x�ٚ�-Lʷ�U̵���jf̬�E��-��T���$��4��s�32M^l1A���:��;X �ys�9GX�bE�]r�N������| lA=��s��_��g6�B��C��^��¡��G���.�2i���ri=�Ve�@v��?mX���S=gG1m!���<�d�2̬�O���?K(�xb_�"A�^ZB�f���K�v����+2�"E?Hyv{����DH�=V��K6�=������|ӆ�z6���1N��{�}Zk�������|����m99��e��������$6@.��)�Do�{�M�"��k/M?��-� ��x l��v�$��f1�f��>�Qu�6,p��M�r���~K�9+Nۭ�D��a3��7V#N�
p;nFK��T�q�PE'4�K��ǘ����=�7e?��T�����8K�����pd��$�kBq�L�K�hޭ}��:pk��@�7 �5���kd:���s7��\�(����}�aʠ�B3Ÿ�C�:�z��tou�8�\�����c�K�*���ęA�t�$�U�2F���+�r��x�guvC���v~�����Ą1����O�b<֩7�A_�%d�TS�#\� .��7��@�n��:b뽷ş�	r�O�"M�0; �W���~<L�!޲Y��<�[���x��F8a��,����
� ��R$���a�3�<C����,�!�BzKز����.e
��3z"rE��M㛝*���bUֻ]�N5�b�*��V�}�>���Z��KB��W��#�k�Kσ�I�J�*~�����r�pu�/�<����}�1{D����6��̀�<�|'�+���ᾐ�����tڍ���[��&��1L����Pw��p}9w6�52�d����<e���\�C®����>|ʃRD��/;��4�8����ڶ3]��l������a��"�%��T�H2xȋ�`p��U�����%6j�"d|r�d!�@?��.�7@�O� �G�9xB�,�o��kc"�~�6*o���l*���A;�21�[ɬ��J�,���m��ω��y���5�8э^�#
=.?u�iKip_�3�jIk���㝿[�)�����u( -86p/��|������~�V��kf-���U�3�+^�5���mx6F����3ᛮ��3(�ߟ�X���И7��4�-P]�!172�	��Z0q��T�ڐ3����ɰՊ���#�Ȟ�F�Q�ж�q�f��#�GÀ�)gܕ�i *T�#��o��}6E�z����Mk��X1(���y_�I!��W6��F������6�9�����;fM_�I�,�yυ��=�u�.k-��4���u�8L��?��P�ZJ܆�Y�]�혌xQ�Jk�/$� حyV��i<*qn8�U?&N�-�� |�4ǥ ��k����s��X+�M�#����c�����l��7u�VuX��NM����iyވ���6��/ɺ(x���#�o���C9*�X��T������5$��%�3���R;d������#DЖ����7�C�l�N5�E� J����Sb�:Q/ o�y1FzU��l�&:����-��2�,��W�#�������\x*N�*�j`�V$�Jn7�;�*�0�+�������	���<&�Ez�Dm��:���At������Ӛ�Q�Y��ŢA2���� �L��i6��W ������2`)�o^?&��~���g��,�ap[�j��d�8���t�#LW���&�I�=r��F���B�e�t��e��+��$��5KŻ>"����ԗ5;��\.����6��I�i��*��v�^���G�6� C�sF���Q�y
ӕ���!���YZE�׺@p�g��D��A@{<�7?X`�?.&"���%:�G���3r�'��C� .著̆b����5��M@p�
��iJ�N�xE"c�jp��a��b��>]aP�V`-��uQ*����-"~O
��Ph�dr=��G.3���K��=eA���P�ȧJ��.�[�O��� >��9�NB5iO�*�^؋@K��G�=22�l鋖�g���|�k�q���jO��:S�!�v���<d7��MM�Wm&ݟ6�Y�����h�)W:�<O�K��o4��>	~��k�����Q\w�>����<�3���c�d�ԸJc�~�-������������
�t���Nx)BX���q�ژ�ꁯ�K&u��/"0��Ge~�F~,\`yTb7c<[d֗�{�[�g_��:����7�s3��}�]�O,r|��;M#^P3B��e�Gi��.<V��a�߿BD��ze-<Oy<�(;36�)p%T6���=�r����o �ʜ�D.�����9���tN��+L�Uw�J�T�S���x���:��wp���w�3y�B�8��Oe���H�xmq��F�Y��tU۳�MN�BBȆuFw�����������/���<�Hy9X㽁�����v�,�M�k&ptxf�nA_�p'^���o�x�l���}�����xU���2I+ЃJ^�:T�~��8�2Ʀ� r�r����	 �i�PNw�$�AiB��jst~�2�2B��`���4Þ�悎� =t���׵���'�� -�g�!oM|�MT����G�A��<g��R�z�ˉqp�� ��U��ʠ���W�j�*X/r�j�בZ�� |9���k�{��$D��L?�lK[��ck������SŬ�E)��6�_8ذ`F�
i����C�d�r����E���h/]�x�N�iMo=*X�lH�����m���iv�'��>��;�yg8k�-G��[�g2��O�qt�P��6��Ц[(b��Ŝ�#y��B6|_��j1y��8�G۽b��Jxw�_�;� ��0�<���^�t:��D�7�{��"�|Z9�D7�.��#�{W-����o�f�1��Ӛ9��cr�$NN�$]�_�s
��̥�v;��r?�h'*���|�9��)Ax?�7��X$�R �sk�;�Ԋ�j��+hu&şfe��]C9�M��-AYk�^E��mBJ��>������A��R��㮶���<���I7��C����a��{����q�њ����2#lYܳ.�G(�Ý���h��l�Cf}���:��Ԉp�F�?W4�Z펾NT��
�eۜ%�Z�s|0"�ae��I@r�dg W��뚫V@�P���Q���~��lP]}ڣ<���ն|]RX��&��a:�u������ě����Qr*@��7'��k��;h*��W��ą:�(�4E���x0����{���y�b���oEP��L�"��l,�T�M���K��}��<C���$F�O6���PU���2��;UP�5��k.4�"�U&�
���qtsS�T��$H��A��w���۫@�ӳ��h4�*?���-_�z��K�@pU�nOQ�ad����wU�����	F�\���"�e��Ҝ��d�� Ͳ(q���lؼ���><,FN��e��	���̓�M�Η	,[��o��j�5����������Z5�0��=*��7	
�d��綑�-�Jn9F	c��>�|���2���z!���	�s�RdT��!0U�d��.�T/��	���x�bۉ�P41�\{jj��0�~�?O�����U�,01�&�L�}���d�n��RE�i��.�k;a��5�V��PGٮ}�m=���w�]+�>���A��h��vyZL�������Z@9�ʭ�D����^�[�9
��`���*��1�˲�G�1�I���H@j�N��2��`��Glm-vP��3#u�7�L��6aM�^5��Y^��3{��L�2�L��j����y0�l|Z_�N�v�1[d��́	���ي��kb���	�����s>�w�@�h�ޑ����ni.I�D�S:Ym��]�~�b3_�Uuy�uf��a��+}��=��M���}E\�E�%b�p��o_��a�|���=>TC��K�<qS(��qw�+��}&OM�C��K��j�:�O='��� v����?h�g:,Z7W��`�0|�%˶s�o�"�+��
@ ���E�ں�M,�?�K��T!��_�|"!�}�M����y/�v�f)�{Y�1�w3�a�ka��\+`J=];[	B�Vd0�ڿ�4������u���sQ�	��#�@�_!�����2R]�"�7s��͂��
k���N��j�A�c���A�l谴D�*�r���=���;Xj�U��c)��C�#�����D1}��PLt&~�IV�~8-l�¬+��Zvx-��Y��.���y�����޹&��B]�\�x�~�G� �y�+��;#؄�ą���o9���>$��4["��mD6�׮�3[^�ƾ���V����v7�l����̠�t��#z	PW(b�Ȧ�_i,�a�87u�� ��{��?����[�e�d�O�HA�cn��qN-�6���@��Y�l�&viM2��E΂)o���n8��
aHg�������6�&�dp��:HRnv�VF^y:Λ-	�;͞�T|�f4{�,��W���M�����	�ɹ��X�W�&�5���T��"��,L�X	s_�����V�	<��U��pj8?�u�	��w�LzPt8��C��xBP�M�2�Ҫ/@��#��F�9xʽ(X���iM�m~��c/��S)�����3�f��w-b�[��r�`��OS0T8�����KT�������#�����c�Xuh�����!5څK�m�rN��D�uȮR:��H5�9e=�����:Zf��aѵ���c�p_u}��\�f��n2��FHt�;��Da�ێ�}p�_�k�M��MF�҅u�OɃ�� II��JLgc�-�q����v=��+�h�j8�����7�]���zZ��ٯ��*�$#U�JdLz�J�G��ӗ��i�ZO@�H@����nX�j�L�Y�k�ʙ���>�ݶo�9`���x/D8xTr��ָ����=��x��� �i�9UլƉՉ��w$-d3i�~]�H)\���Jѳ��߆Zɦ�Y�`�# ��ÉO�wY��K\Gfg+?ʌG%��Jwy:~�Ȃ pgAlSCn����!C��Y�J6��d.k�7����u�A?�"�"y\�Y���Ll�\yb�k�Ӣ#Ys�Pߑn0�NN�����PxGg�߫I>S�HQB�v�U�;c��N����A+Xt�ֻX5�,���ê�~�o5�l{�����匒�|S���~H]����o�8�������@'��`�&g/�`�'i����1Q�;�}^��پV����<VwZ����>�C�\�o����s3�"�%��(AxM������n���=�����K��c���(�4"�y�5��ŝ/�)tՌ�`�>C��b�]p��¤�pޞo��W����VYJe���؟�G�"Y\RM��H[���P2�(c���T�0��E��*	��g<wb];�}�b4,��@�=lsn�3�?Ek
�rlN<*@£Q��F�~��On?Dt��c�J#L�i�\�5�>r��׌��'��M+�l��P��5)ʄ:�����sj���j�9���b�ʂ��Xk:��6�AY��,�~��g�gR�5�XƼ�:fh�O~8��
&�GqK"Q��8l�ܶ����&�`����ܸﾐqm��kU�������\�٥a��<\9���t���a�~���V�i���'u�4������d�e[���<Av�8�5����9����T�Q��
 p-~�`+^�\P�S��8Bd�u�+SO��KR�F�}��V�2�]���ԉ�����8a��p��ftz#�o/��ǮRX@�����4�{FᢋbxU=Կ��:Ӄ�d�'�c�?��Us'�s�|�Q]^Y�U���?�>2t�6��e\*ٞ�!��+O�i��{�$:�{�T
�΃�1T��DE:�7��F�-	y��3����"�<���9}D���d��0���9(c���e���4��,O_��/��NL��x/�{���tۭ�0GӝJ�k���`{e_��No��P��rD-,��g"��8��,
I75Z��
��5Q�����R� {q䫱��<^8$l��&,��s?�5�r����/�ڦ�Wo3�-�ހ�T���K��`�'�!��F֕�!I�D����t(��	��%A�[�[�>3_�?۰zTcN'��s/q4�D˿�X��ܰ�7��[��?�N�8)����
j��w?����H���~9�O/�[QU~w�����0���$��i���Q���9�E��o�."}��@aSo�U�{y�6h�)jJ��,�u%9�cڿ�������f&t�2YC�)[Њ�:�Ⰼՠ�����2^/�x̡��b���q(��	/3����_|��L����R�����v�F%.9_��+g,�� ����A��M������	J������6=rE��e9q���~����&
�;h���N�T�ʷ��C��1��	+X����I�y�9�/h!��p�[�d(֫��ڹ���9�/g�f��Lt�b���|��?��=�NK֖h�e�cs�y�;�(UA�������b�>���8��s�Zl�A�Xb��N��_�K��t��h�(�����6E!<�\�����z��-�Ê���fna��[n@q���ٜhC���^h�K����(�$���p*3�na٣	��p��f�<�W��9�44d�(�#�jN�~a[�`K�E����K��nrr�9�����I��o+i�:��kEcN��|�%�/|����)���e�ޜ�eŷBR.����#P(dg���P�:��hGe1m��/��\��ݥ���z�E��0Ek�A�\���݂���YZ�"Mesk;/��uNlF��c��w?N�� �v��V�R�*�v�����8���ڊl�����cXpM�Z�x�_6�2�eX���m��a���d��(�{�a;�>�I]j���bw�;H�8k.�M_w�kv�;ǭHW��.&t�ߡ�<J;�k�%�����H�D���U�m������{Q?�.O���S�Ǎ�Ak�1#�^wʹ�ˑ
)�q��5l��ZÔ��l%��_E��w7ځ�Jz8�TL?-�o���ğ�K`�ԛy�(� )*�e�L��0,5�.��$TG�9$s�+�"�c58솆��ԇ��о��/n�J���F��E��� �'�p�U��Ȱ�T7��\0�8�;��G���R��.k�%� ��O��I� ���'���C���p?���1e���V��f��{W��O§�!Xs(A��C��'�)=�l��qn���3�Y^t��6ZH۟y��N�C:�UO���%�tU�6�$ u2�)����z�/���T�K���Ȭ�R���-�D�i|6�(9��F�������4;h�+C���@J����H{��ǹ���Φ����:��$@M�֖�����(Ҩ�W� �)c�>��̭��O߅
������4̴��3,m��bq�L ;�Ӭ�t�2�Buv�	#���Lq��Ȝ��fd���7M���!hX#q.�&�%��_���∼�Q���pu��y�r;?����(��6p���]�Du�G0����L{0��`&����ECӌ��nz˷��$V��(pe'Dގ,���H�B�
Q��}TvsfJ¥�<UDQ��:[h����UF�n�/���s��t�
6	���)�������w��-�X5���Q�����1����l� $&/�u}��>g�1���t�	�*�YQc^��X>X��4(�W�|��'�h{-�wj�m���f�O�*G���P�g�͔�ӭx%�l7*�-��iݭW����	���궕�]<9�f��FpoQ�ȶ����y�.{�x�����7�ݫ	q����u���H��Q�-��}��V���BPs���E�Ώ������O���ѣb��j�@u����3�����*<���3���AG��k�=�^Z=C`���8�.������ï����:���x<&���TZ�M�ȓ`�oXd &�r�}MR�^RU�oa3z�f?�g�r� *�J}�����#z�d	��?�e�c����	�L.�c��d���UEѤ�X%�|'�G�%w�?�U�8��.�1�"��vƋl6�m뼿/��z㥢h�}F�<���#t[C.centͥ5�����o�H�rꂵ��s̎4/��AF(uG�����&��Sh����0�L�5�k�<�B��~� ��C�6ݓP���a����${�g;��p�K�z�@�:��Ѐ�5|�񹊭ΞVK�x��B>����Z�@�R�{�C�2Y�c�R2ߣ}8�A���7����?�Ц�ʚ���PB�%�z������/� 	�5Wvx�+����v�?��ș�Ku�b�\gd��
��p�MFv����
8�pAj�ѓ�_�.L�l�x6����V�S��h�.dGbW�T���t<��<�\Pd+0K?��d�Ҧ��������4µ�]�F�>^�p+����Q\��� 2C�&-��xWM��؋7HLԁ|J;I����єH���dg��G�^^�����R#�o�5�l���DH�F�zҡ=7��~ei�x;WPZ
+��^֫��U���ZE['�5�5�����������s��ԃ �������DUQ��
����r�����[�d�k����7���ZB�	���U�lEyp5#�n;�	%\�|��z;z#����z)ݭ�rک���I��Uam �Z�������R���#g��N2��8�H^lP3�Ju�[���k�g�t��{Ѱ�@�J���1)C��߽�M�&�?{2�*ۍ"Ǒ��� Y,޶e����&er��:EV.G��(=mYE|���V[����6�����_���͍��V5�nlNO�>�Id��̶���Ũ���斺eCB����|��-�#(�/��hц"F�Sg�?ƭ oYՇ#+���ח�h�5��S�O�A#�t���o4���e\�=�x0�Ba<y����Յ�	T���%s�h��	�)�hn����m�8���$�s�K�z/�J2v4���#K/�UiJ!���??��z���j%� g�g��P#����^�,ج�\b�M[
�y��<�$eQ���ؖC�t��9�oWtUW�о/
^�+����ʶ���B���@n1w��<�h��DÚ�CY�T�2v�2��skuF#���`����*��p*r��=7d���� 5w�� �
��
!u��;~s_%�;�N�~"�|�xD����$aG�uz9�����pn�׷��m��	�����}}��O|l���{�V�WQ\��u� $2�,��^��`�L%�7 c/�P�:�Y6��p�]f��ZRS
(�����x�� ;h�-�lA{('A�������!��s"��+�m�9<ӹV'������n@c��m'����%�����FZ"�z�H\�<�}��E�b�"N'q�43S\�Ѓ<�d�ig+�Өq�D���4��  <tƺ�j��c�Ņ&M��8w�u���`K`��%A'B� ³sO̬ym�tN�˃f�mx�}x3od��������'7�A�
��Rק�`�'�L���3z��ǚ�ݞ�t' J{qZa�n�VC�V�c���n�+m
n��?�>y��g�8N����U����4*:�RS�n�=�&iM���G�1�p i{�
{b*�̆Y���g��d��K#��v���6l��Y�,>!�H�|��tƛ��%��J	��p��ҕ�5탹�F^����]3G��N!��
�D���ž�/��}sr[s�e�=�T�h�������d/4JZ���c���Pg��	���?�q��wLf�h�)��[Qn\�S�h@�Y������w�4�1�G��_����Ƕ���:І�F��������8�Y���;*�{�����c+q
�]9Ȑ�����p�3`$?#���^��,�^���Ǵ;���F�2��m
����o��Ǝ^p�57�H��i����*]�l����r$?�����lKO\�Az��uc�]4�)��o`*���$�������f[���ݙ��I�eR߭y|l���^�����*jy]�ݔ�j��7P���.^Ȫ��{~�z��L-�Jf�6	o�fE�u�Ӌ���H��[8�Hj�o�8����{dl�|���a�v)�T; An�lɸ�=��)�O�⍍�S o��T��н|�~�6jLz1�-$�
��%d����K�� �ڵ��'��ak�4����rO��Z�f��b{zFU��ϵ�?�cc��܎��Z0��r�������mo_3۩&���+r�����y�[�����b��#(>C��<�� �������i)V��X�8`���н`7����z8!]�s�T.��H�����n�p3qR
���}�Z=lT��c�~_�8���Q��Cȇ�S�����Vji#E�cP����o�&���K�@�ܝӫ��^"�H�D��G���V
~�`^�G(l���)�(�d�����|�ٺ�S�b�/��m�Ґ�B{��U�P�=Oo�\�W��>��H�
�N��G��@�!@���_W��D\�~AU��iא�cf�e$����Ը9���ZZ.��η�z*�����z��M��� ��c����&��/)��<��(k,��x�� ���Rd�)�lU��E)�ׇ�9�"i$�z5ۛDlx�S�5��(S����gM	d)���0�x��b�|4���>-!S�)�a���+?�j��\�����A�?KY���O>��������tŋsw�ڬ�i�] ��AfY����sK�碊kMx�±���n����%�?����e�j?M��g~nH�ﾲ7�4Ys��͏�r"�\#�
�]^��XY!�}��]���p�r%j�MZ{��9��!h�9<�4h��m�� �������\,b��l-��mW��j��-�h��N���隘�	�>t��t�9��}mޠF}���PpӰW��'�K5~5�l"����U���$Tm8��/��P�dC|��[���Qx�"77�A���v�6��z%<�"�`��,� [�\������>x���٩	I��.D��6\̰�׺*�\T����D.��@�	g ����7G��%� ��m�V�q�]m!r�J�k��\��F��gI��)K<eI8�"[D+��L1������J|�ۥm�3쟿S$~@3�PR�P(]ь�!�{ob]���fR�q�׎#�i-��v��wc���u���@ ���I©�����;Gd���%<V�o8d!K
�����M�
�ΐ����P�`�ѕ0:}�<�U�vm&@��+ v�ܼH�L������݃~��k�lks�J���d���)�\�G��l0�f��֩?�0�C�O%mP��3��;-."Z��ctD&�C4on-��lrL��X�!��l���z�o�X��ٲ)(�0*�9�$����/���9)N�A��"Cʌ��W�q���,��������4g���P�PtS��]SC����̨��Wh�{L���4�)�Xb�>SC��P�)Q�X�G��L�@�$�<aų�.�|�$�������W[�&�o��'.�V���M�uH�gヴ!ӹ}V�"?��`� ��ʙ�Y@�9;Bn x��I������1�\��V�H�I�ڀ�������n��s�����!
�	0w~\ۂ�V�;�^�sxp���Y�epb�:�v�E�+Da��׮�2�=�$E�-r<�~�@�Fb�&�Jy~�~x�'�u����7h��kA� �,��9F�l�}�e�1-��D��'9Q|�_���C�	硍|ԏ��@c�G�������LZ��/��h�C�Unr���S�޴���)
2�P���l6��C~#	�230��\;�sy�'V*h��,!㗒������ǢdY!���%�y�`�we��ӂ��2�H�8}��.��r�Z�7�"�h����Gp(Nd�V+����.���e>v���"�%m�- DaM�D�&,�$�Y2��zFEjl��R��"����fi�˚�y%�dj� ����qiֱ9� ��}���\���Զ�{f ��AA9��2)�]�+]¿���W�5�R�K����C����AP�P���v])�w0:��-5�L�Ɉ�.h�O3 �-�e�+:t��=Ÿ>-�+o\�9`�g����浴	�O�ы_q�Ykuy��ҡ���y_��X�!�T|��e�F�i�o�8�P8�c�Y`s�㯎<��l�����*�]�Ə�O�y붧��irޓ�_p��U��j�AoV��P��T���u�s
�4�a�-�1�%_���z3��֮T�`��7y��u�8�sM�]�ߊ�i#o�E���m=9�۵l�,�~2�\��
�g91�T���5������`o��,�I�e(x��O�L�w��k�CT�O1]���5+F)��ΚW��8� @u���P�46x�"�&O)��`��9�R�ߪT�Y� ��Bn5צc'Ie�\�d=�� GpLP�J���V�^���U������[��y��^���$�_�
!�fSv�&XO�����Z[�ܲ�����w��{I��n7����C��X8^K{{�ɊTBxs��H܁	��O&�G���Ǹ�Ap�B��� $�h�]Ur��"p����ma��r�5{c��)�D[�+Զ�D�S�R`�naH\N_q�THPF��If���f]�@��gj�.����� ��1b�1iK\[ӏ.ǽ)�#��i�@׬ܾ�m*�u&�Pg)����]��n+�)�d�i����@��yg�eR�<]L�c�z�Z�y���[��[O-�qd��dra��(���1+��97�3��RS�Sє��(�ξ���m	�l������awZ�S�sq�YC@���kaH��Q�vg.�5�+���~\�� �F	����r��{�8�LK�b�����w5 �
��Q0?i)5��w�X(sZ��E�%�s��� ��z4��RjM?�&����A�-v>���V����#�,6����5[�h��=��e=K�-�ԡ�t�.����wOG9�
e.cw���e}����<V�c����"���gnؾToA���2\��FK�e�'���pӨ9W�ԥ(F�!D7g�ׄ��#��(B�ef�Y�ߑ�,Hr�@���J�0ZS9h�S�<ya�qf96��j���n7��7J#sMu�]и3�="�Y�i7�S���{��X^�
iXxU>3j�����	�m�z~���ܧ�Rъl��1qT��A��Ĉhy�/j���0�đdŹ|��"���L�U�k���r��aI{M�U��hG�P�5�Uk���`T[C��a��@�|=��S��^[bu\�x��i���:?�o-5C��Zȧc�	����fY�T֏�(c����ҩ�����r�5��Y��bh��KY�ހ��ڒtR���NÛUFE�P�9>`6���e�����W���#RJ|\*�֢�+��I�+���~H<,��	 0���ofR)�"L0�g����6f5kw�D��L�V]+�=����T~n�i�<�n��:enZ�( �)�}}I�*�S~T�[�:����x��qb�~w�K�����=D�mT!3���3���^Oug<�)��s�<�db}փ�tGMi���3 �qM�=B'.����\�.2xQ�γ)e2��|0����!�E�Z� �s�}e|�!-�-[��ln�'�P�z�J0Y�M9#q�oۢU��°�Ā�o�2����K-)+�����ę��K�m�ӹC������g��C�׬��܈N�S�\��|�+wrK��TD���`���F�qo*;u�ᙇ�S�L�r�2�wrB��I|s�#cM�˝�iy�t|S�5[7 ��Υ�z��T�r�Ħ���:"�vk�$�:���P%gH'�c�]p���ua��J!�O�H�Z�ː�&�1�ܡ�2��z�Z������X~�oi�u������9c�Z4�� w�,�U<�g.��A�@��+|%^)�2y�O�>տ9���{��̹P��:��zxl�,���iQNt�ta�=�0��Q$>� �p�&6y�\*s�:���6�mH�'��o:�_���s�sP�5,�B|��?�χ���,�g��F��zWM�';�3�V2��5T�vo��Y����c�{��XƋ�2��s!���#��F���+�z��v	<4|W�u���&$8dr�}���\��$v����M��h/B�L�S�]��k��i�ѼU<a���C�e5��%���:�X���6�����/6�O���y�[����&E��9�V �&Q�����@S�{�v�(��8�<�wܘ5��{��D�I���ǌN�x_y%{p�(=�<�$	%��r^���t�`�L���et��>X���T�Ŋ�"J�|jvV*�RDCZ�}��U�@���m��Ǟp�Γ]+�J���)*ݕ#Ef���o.�cN��ǔ�����(�8O��j�}�֤b/���e���WWq��M[�^j s2�8��"A����Y�8�]���
��ޠ�=ۏ/�d5��a	����w3:���ϓ�P�cj"���w�3�睦�B�;A��Ӎ��Y�F��L��v��jP�.�l����OG� uڴ�~�yC���`��dX�]���0̐m�L}��B��[i�ׂef��K��h�_x2��1�>�� �F$e��kU"y~"�P�M�5ѸN��uq���ܩx'C�(������Qpt?������~�*t�|���)�)b��[�W��F��>ҡWB���h8��{Z|⚖l�ãcΉg_���qxp�����WY��QЁ|pmr����K/Ӣ�V��8��J�� �2�ǋ�A-��;Y���|}f�����c�0]i��H���㓙]:䒘�����gʶ	V�K"y�%7�ɚ���z!��x3w~�5"{;���q5�%2@9wR5?=�0�:�u3)��;��P��vc�fw�t塎(QiAgm|��;��\����Β�T0m�w�NΣ��㛩���\Z݂'�	P�Ȯz�0�	��WQ�B�﷡BFۅ_�]~����|�moq ���U�� R���3|I��X#�k6W�G��>�s]wiq��>7�QI�h�9��%�Â�EUI4�<V��CN-=_��;g~`S�w�3J53��1���y?W�#�l$D΍�:�G�u�X�G��{�zC���������!s��m��A����JM}&)���P��F�b50#0��]0[P΃0P~�D��㸕�z]�tO���w�d>ؼ?���+N�V�]-�By7���_Ƈ��&p;ɲ��*��\X�]o�e2�s7`�	��+<K
��Q�`�7��0��ġ}	��8�	i�m��xX�/���U"�2f<�� $�"=f׆�3�ا�)C�7E�m�a^�CI���:��k����ۀ}ʦ8���>���T�7f�9:.!0Ե,>��j����gkv�o�>��!�R�6�3�L�\��À�@\���Q������#|���N��tc��U���NN
%U5��5�.�d^Z �-�Y(�w�$�6�bJm<d�O���gXP�z��O7
H9�YNY`.Ac���Q��T�]E�2e��Օ|����uz�nI�On��A�KM�=��r�;D{��,��فY	�Y�=��v��0�+��<��o(Q���q��͔3�g�\�=�;`�IS�2�N2/]z֒�����t�V���y��l�J���1N_ -\Y4�����Ϙ�M?���۔�É	v�µ���$+f{�215�a�'ab��+%
ԅ�[���46Te�^�7F�=ԭ6�wq�Τ4����":��w���W���qX�����^w���.a���m
���j���5�ɢ��0.6��c$� �8�[�RJ�YǪc�A{9%��%�u���[�|�V��Oj�i
B��%i�͎�o�<��A��� �u�6m�n0��8E�����)����lg%��K��MNA���GO�/��EW��L�Ű!���	G@�o-��.�\u��'Y�V�%g$aP��S7����+-�^�w��G��ڦ}�����Z�A*<�3�NBg-q�c4�D�Q����j�ٮ�2zn	�fM2�.�ҙF����Mk�{��I'��Q8$|���W��+i�ˇV�zỴz@lOb#z�%�փ3&�T���48�Ib~dECI��6�ͩ&=-���L��r��y5��o�N����%J׆VG$$2�K�ev'!3J��	���*~�����z�ә����G�M":}b�$����d��O�wn�R��OU2��޳�pL�������n�1Hj�Pu�6:]睾�~9�kq�8��l0:��MWE$|RJ��\f�8�C�����(�vۇ�V�<ۋ�h^|Z�Vk�ZòFP��G��Ƴ���`��G�'Cu���8K%�T�4A��;��,� ��V�Ae�:Z�������k5��@Z1E��-�� F��Z��aX�ӕcK��Kl�K��
 ���P#S�R�>���z��FR�&֪��Lγ5��� W(C�>�: �^%^�٤�M}���Mo��V���Qo�Wh..�T(>�Ĩ4������'��<W�u	�qHڴ�:*����h�\��mJ+��8�C����*�5�'u��E�Ld׺��	��kF�^1�R��:��Lx'-R;	��{e[�FXe�daW0�����d���*��8�zUw�̫�R�n��"Qv�0�ԫ
�]q:_WR_- �vb�+T�+Bz�ic+L��&��2�D�����L��%z��=^�L���� ��Yq���?B8�d� 7[Bs�R���*��n�op�A�Z��	��ぴ���y~j5eW�&���47k��?��+>�]p%�Ӭ/��
����&1�����g���{+�M&N�\:�~��C ��1<��>!�*/�Tm$d�̀��bȜ$��-}���J�:�mK�6���\о�p�d`�¦[`_%ܺ'n�R��p΀�}�b�"���jː�����=ߎ�T^ R��>�_']`(�>�u�R^����3�r��4,��X
���޷��fl�j�`mu���ͬ��-@�4���#�O�kc�g�4�xS�%h[G��!蹁T��<���Wl��%)N�1����7^���r��{��0�t%��
��F&<⢜�2��O��
Z7�V0����a	�q�V'F���)Z<ڑi����Q8~��k�NE8Q1��X�����T*D�ӯ�BPi�'��m��ѕ�Fz�|{��x�6@�!
t�#���!ܚ+��(����:S���%hJ�f����/ ��l�PH�X��x���L%K@��!A�wx竈��`�I(�DO���ք�'q*����V�(^˃����i�\�>w�2�]t�ؓw��ߘ|{���NsO�3n��V3������o��9��_b��Z7�z��!`f!5�2�N��6�Ɋ���<�|�D`J�FH#�p)j��LP�I�6����X������E� ����5����6��q:����:��W���q�xT��sQw�������<���[CNcw��W�YB{�{$ܰ�;+����72����M=�ʺdK����M�2�٠�疲��K�lV^ک��VؖC�z0��A�!3X��[��U���j+�+����uy�Z���4�7
�+r�J��Ē)OgR�q����q���"�A�xjp��a�Ksv�
���;E�!����Ul2����YF�]_ٹ��Q$3���t�������8ğ`�������2��姓CY׼=�t�նg!�1�&-4�1��ع�C�z��z���N������+UZ�[C��n\�v����tHK�t��[�r~b2�[�E��ǰ�� �*
o���
y�4�?�����[��	M���������ծJ]�ݴ���bfn^s�Z���d�+��L����%�'��h�߿N�-Ő�`=������-��2�(yq�C�`�+���oe���6�,.u����!�&_��˧�^�[���8xErS�h9Ղ��JyTu_��{�N��k�
ߎ����:_������iuI�YF���lyw��fF���&�)�3^E�{˃��<!(OO���V˅ ?HZ���u݄��"��urϗ���]��r�=��@;��H�Bwކ��y����`�,v}�Y�&A��~p;�.,�k(�E�nzєMI��F(�v�+�N% e��`��_F,����9���(��j��/7�ߨ1�r��g����6 �[T�cO���l�8�>�e�bmÉh���� <���ǋdF3r+J@�8}�״�rz��t�Ԥ�m�l蠁��9�
;������\o���m�;04V5��3�ܲ�I�����,�*q9h���0f�ol[���iv1)k�lo�.��CL����Q���G�d��o�,�L#���)����yS�c]4��(��LЦ�a8lt"��1��,����{����x��O&��p쇓����?��OQ�s=��`�#ڲ=�C	��nB�/K,z<X���5kk%��Az�H�6�0��셀I:/�K��P������	4$���GT�p��T��Y4MYڼR,�(%���Ĩ3QF`(MM�&:qȌ�Q��Ѡ\:m`��r���QU��d6;�
?��^K�h�W���}��JCf�a4' �3�ˈ�9RMw�����ײ������+��xU ��T%�Y���e/fh쩿"A��}�mJx~mxj5O��Y%�}��FU��������٠�����!������`S�R����7�i�8E���!�?���h$�������}W��9���>�y2�#�6�Z&����n��{kuC�`L��ȏ��}����tB�?�up���φ�z��W�����qAl�bH���I�$i�{�y����r���FC�a@��>6 �ѫ8$ٝ�<6���
8��9��5�I�����l��zq�3�ڼ������z6���F�#A�Aa]�v�2��%X��w�ť�Ղ?Œ�$\$0�������0A�����5��
��J��܏���w�v=��΅�~sw#�oұY��M���-��o��ጳ�����U$ŀ��8��D<n���[*Z�m��T�g��j3�����>�s#"f���PW�h��^�����Z\���p�=�dM�\"'��q�y�w�95�*<4��h��u�+q�S��5)�k�y�Z9�N+$�r��dc&�g�A�]������<�������fJ�|�eu�@w��z�.3��Q�&.����gg�����%��o���@'�q�5L���9��ƢV��¦zR�_�b#*�6`�3���<G�F*��[�܎����Y�s�_�1̧m�M�7���Z���㪚�`�{c�$�ݏ|�|u�V17����F-�hDA-��Y8���G/i�c��x���	m���߁��� ��cn"���L?Y�J.z�X�<�
��5�9�|9p����J��������|��PZ�7�69%b�DJ��ߥ�Q�6���\�J�fɡK~_˓Iq���TH<�i7������ź~��9iŗ �tk�ۇu�%�Ʋ�$�p��\RC�S�l):����񨑌�F=_�Օd��2?�T��� �����#�w*�Q��m������,��
�m-�߱/���abh��S���v4����?\��0��m���X=V<�F�:��&:�,�"ڔg5�%g�% ܧcjd$'��r� {m�Č�� /���qz�
�������ɇ��,Zu����Kh*�!�<�[��w �^ɼ�֪�V+k@�P�����zG�K�{{֢wU&Ani[u�S2#���������NOK������¼<.z�3� 3'O�yS�4�P�a��nEX@/�_ >3ŝ�к����P�#0c�S/�˙׹�<ÏB������%߁����R:/�4}�<8�����ˮ��ӰF��2��HH��pA�uױ��ǖ7�s%�����Vx��߁�e�a|"�y`����Z��#S���>s���}������[�ӧR�t�Y����w|���q�Dθ|zY
�7
yy്xZ��F{����>"	��W��P�}hˇp�|x�bi8�84|(Y��$u-�v�J$���Y����b��-S|�>��+?�҃)Q���U�F�Tg�ݦ��^(��<�jA8(���\�I��=R"�B�y�xp��<����*�T����t+�*[/�c��~7 Տ>.�X&�0�p��I��P�==�8c�y@06善�>��i;��a��<¶�^���R�[K��.n(���>8������tl�u#�c0t6��b�B��)��볔�*U�cc���]�ȇz[۪���GГb�F&�t�L�-�w>�/co6L�?^�M�T��~m�Mf��`���=	�~�ZD�U6�����4���맪����H\TO�c2
L�q�)~C�xǿb'!k��p�wV���JM��C8�~�:"U��;��U�9�.ƥ�	�/��4;��'��$s0��J�ρ�C�A;��L��s�v��PYf(쒈�W�l��]�*�&�K{�;��b��)]�Q:{�(S���۔��!�߄�z�ڀD�� �	��G���a���&�h^���g�?�ۋ�*8(a4�cI��3*�f��֪��7@qj��I܅.�q:&��hGAcUv�%�s�uI�㵡>��!����Q�J)��)� �����"G��yW	�H��\�k�D}މH��8�{$�k��a��CZ�0�Pc�[���s-�xv�(��U���2��P�7!?��[I��ЬC�:*����˦���RSї<�M.x�L�ٰm���a��A=�S+:&�x����U���z%��֦%�����t)_��[��餐3��q�Ϣ�Ҫ�X4fc�~��p�I�tqcV�Z��l��p�ޯF��g#�\� ��/ �r+U�<�9�Ѣeb�� �J�+JE���>��Y����4/UK�u�^t`B����p/׵N�n,�K�3Mj��,R�R�`P&�%�x�FɗGI�_��}4�3d�DEt$��V]9���S%u}+����'á���7�0��0���L��ܔ�z?rRΞ5�L�I������V[��Do��r��z��~jq�a�>U���]�fIn@�����9
#�.~Lh��g �R򆮵Ź��L8�������c�7%�@s�PP.�^����.)my�R�j�6�Mj�!���#U���sWP�A��S8y���.5ܻnC&S����r�
�����P�����?*�'^c<p��ǖ� Kg�Yt��|�r&�O�0U��~��O��i+��Pt_��<Z�?�h�E��_�v����@�eR[*�����%)GՐ(kS��B��Jhf��W������"�<f1�f���L��}�D�|���M)g[��N^��Rj��W�#4����SC+�Xn<k\J��*ڨ��CdԞ�*U%[�����)����0!��.& ��JZ�:�=u�'��ݹ|�oﱢ��;�7�wh��40�o�}�9|ˈՀ��[qPT����L�q��(k@9���*{Q��h�	=	�����q�0�/�zȄal���p.��-���r���){C)_Ȥ��Z��cC�p�c�(!�rġ�;
W��@��g~ވy!��������;��,�#Y)]B��~���W.����x�Ɗ�)���U��x��io$��3��Z�JL� ����hg�����E|���vK������p�K)mZ��P p�!�q��h>�M��U�4�%R��*a0���_�1�����(a���yU��{��T��[���[�Oٛ\�~Z���7a����^H��$6�?�2�aO}�yZ܃7�^*(`	��.�7�!�H|;�(�Ef;$|U����#��Y7b;(��$_s�;ARxG�Up���	���^�'~%«?XK�1����ĮZr4�c�X��W���u=�3T�m�&=�@���#à������Q�H}b��]����Lѝ���"4��V����b�\�_F��p!���/�R��nz���?�h���_#�׹�07 Q3��_�Y�+���J�MO}V�L�>��E��i=��ވ�f�r��t�eo2��Q%n{~��[ܟb����2���^Guk�H���=�0����7��4�`wr�?�>೚Ke�-�	�IzU�QJ�L`]��W\���-�]0:�RB[�$�k. 
S����k��
I&Q��g��L%��][�r64��sVm�K��E%�K�z�>�%J�����TsK׎�զR�d��Su�����E�������
�N;�Dȍ8�1�'�F�3��yP��I���$�q~�����l�\%c��4���	�l�9s_��XI�e�L�~t�Y6<8��Cާ�H̊�b�X�c@���1,�"�<����g��Y'b3|�7��H���3`�+G�=b���^�K
B)�>#U?"e��C��c��F�ؤ:V���P���M޵�h�sl�{̚����
�jg;�Y�5��'b�O��g�'f�C�~�uD�m�{2^�����$XK؉�7�jR�eb�y�'�{���a�8����D%3��V�6)��u��vᲲ�s���,�
����P����y�Β<�)
;H2��-��M�^x�+�L�+D��WB�,�Ւ�gӥ|A�m8�h][��fy��c�E��<�k�|M5�y�`r�L0���?�񏥮� �d�l��{�a��]4�� ��W\�^��"MhGqT#į��UP�-{[Gmi7�,렄F+��>���!W2�O3�*W�����v׼��K�K]�%b�QU:���t��.���,�����������0�ͺK!$S��ȫ�-�@�:�@��D�:o_@s� 㔪���c6�qrYV����;e$����nY -uN`���U�%>�����	�9�Ĺa3b;�D&�1i���Yt's�M�zU�)a�V"�$�~F���(jw��/�[re�i5�8f�q#��3�T���(=Χ�v��-�7�����<
�f���D<CF�����W�=YF%��V�;�,���ݠn���R���N�m�K��J�������stx�!���BaA�|=���m�SS��%��k��]I�8��Eh1�T�9*kt�g��Lz�X��&s�ܖ�y��D�MC��/⡟��fZ�����E��}�p-r�ժ�by�U�f���&�X|;x�#Qڨ�	MJ����/�H�����/�䲶Y Ï>�}ЁJ��q@0�)�^����k*K�2NI~Y*6�U}��#��H��1���~ ����s�JԆ��f��,ٍ�أ9~˿7�7E�`������,�{��0��:�����7����_Z�\S��I*(^�W1l��2T-;r믩��~b�kÏ���Js���,j�Q���cs���$���ZXY���Qχ��MecW���w�b��nEVx��&��HZ�M_k�6RB�v�}f/��;���I� ����GO�3/<���u"�Kd�"\���m�S��#,��L��I�T�j����_��	k������jf�O�Z���`�,�ޔ����u$K�G]r��'��.�<����v�?%��U*�=��c��@cfXfG�"L9ɱ�����>%�g�����4|9��*"`Z���c���Oh~ h�&�ڹ�̚(v��z��frS���\Qw,��N�]�s�DŊrq9�-5/�*�.�*��s��x�jfS�phH4"u�cǬ�ȼ|c�j8��ͅ�@1ù"
���}e�Jh$9P6�t� +����c����ͣaneS����E�VJ���V>?�m�>��e�(�����m���RB��oo���>��E�Kwb8%RM\a���#�*Gdo�'�� (�t��	@�zl:�ß �����p]��_���굹J���
X<�o��OJ�����7R� r��
L��1�܃e3I&��TK�c�Q_O'�tW��&VO�+�K,i�hz�jl�Lu^4���ap��+F:�ڥ0��ו}ׁ��$�!�����4ʦ�B��龎�PHf����<C���L	��d/�W�Y�wj/����N�3@�}��>'<yMh���J&Ƙ�$�>}����g(ϣ#;�^�����B7��U����n�����l���9\��(�ޔ�?�<Òa�Z��$�a27�$�l��ط^�V��;4b�� �GKK�b>_.s'�#�x�W�F�H=N��Ճ�,nc	�4�%
_�1�=��xM�̼9x[��mz�<	w9����\�q�x�
X��"�	<���9�3�_<,�0��qi�.�b@֢��-�_���K[�ʹ4���,�$` �N�y��?,�����'au�#����OM��o�=Y&�ձ�8���b-��j��=Fh�T�����s���٦zx́|�>�����#��>�{��zc�A�1��F`����a@5�04�y[~��eN\���N��������b�e���s�'vFl�pN�W�J�̼�E�u��̓�S�2pK5T��#�i��U��W��h C���w�}!��_�ߚ��
�֍w̓�S�����3ߒʩ�"jiC#�I�A��2\ ϶Q4��/�����Tr�kA�F�zYM�b^�
�fL��E�K�븚�Q)�07{�xIu����0��Q�W �辏XF~� �a�g���kyz�6�������kS�@DrF:��t��"��-Df[�gs�Н�d���f�ٮ+��U	�[8���%�B�S��������iu�T�O:�&��k4i_���4�{P������{�2���'~�A��Y�q�=6����帺���Y���cwGW�� �s�\zO&�Q�ءu�{��n�B�&�Ho��ji����a���h��E< �I��n��e�.q(+&E�c�O%q��3��$$�u�UW ���R�z��	h�@oY�@��$|
l<����+,yQ��ep�B��s�Ku�[H�]S?��ݢ5����m���j��/����4���Z�Р��C#¦�Z	����U`�#9U�'�}���������u5xU����Ezz��q��#���70]�o�>p٠!�>������C�߭K��h�����U����;%8"�)�Q�n��?�H:����|�.�3o�Ia��Q�^~%U�-��Ѿ�p��I���TW̙��Y�Q)��-.Ό�t8E��?�ݾb�5��p�W�v3�;7R&�]�A�a����$�˘�����&`x8O�Ԏ�m�"F�W"�����I�*4Fm���?B�HA�,�y݀(o� ��眖�*UyR#��k���C����� 0�|3������X=`���l���m��uqH��������4�i��2���,e�}�/O�M#�{�����=	p�Yx��Z��r.w��Jh�`c������{�c��fY���.o�A�#ō���)*��	Zq\ޓY��K0�&�'A��+�H�$���s'A=��!�Ь�}&Zu���7|Y��<��P����/U� 1��B�t�v f�1�2.�3�N؇:Q�nG�r.���j/6�n Vϝc�nm.�̔4�^�\k��2�X�|�{[L�X��AL����F4 쬛'��Y���f���~Xp@�\"�����޼>�ٞ.��!�SJ/]�GQhqQ��5���	;p\Ld���]�ǯ/��v���1��	:���c$�����	�nEҍ@,�����a�l�E��A�0���U�,�����A����VP|�����,�b$���U�װ�j� f��Y�)���G �:u��Ut���
�1Oͨ���!�1��p�(��ڬ�����dZ/�a�"��y�D?$'�G1�����j��
3P!0��7�9��:v!G���X۾9.��[���'ݤ�ځ��`ШݙO�ԐT�aYD���3���f��c�1�]�0��uF��	Bqfԏ�:L��Ȝ�4L��i�_S�i3D��'p+?�����!�٧"R��LS����6<�n��Ҕ�dU�{W�oNB��K�����,��:/Q
?�|Pb��C1����|x���hk ���)����݈7qN����'v����-/1Km�*��1���k�Ԩ:�<j�7��#A=<9a�8��uNh¾�. ��ơ�.����q����"�Q�J����6�
hҹ�n�L���WsbjM_�_�jZ���;[/#����<��۪�\/n&��j�[��ku�Vc�k�X\�������B^��F6�s��3c�K��PX�
o�to@a�c2Ro|������d��2���u���=�,U�t�2ǭZ&;������-�^��ntuc摳���uX�k��X�����^,+Ő��[�<��,���̢��>��cBd�a���5��"Z��)W6"$�q�%0����w>�wu"I�h���Ӓ�?�~�5��Ȝ�=�:��VZ;��Us������� ��]�E�����(Z�'N�m���s�6�6)����G�#l>N�ǹE#0�io�岱��{4y۝j�^0�Q�Nw�H�'Aվ��3U�8�ߺ >���	�,�˷IM������� ~���V5�2��Pe��bsP�t�	u^�����=��xl,\�����pmEZ��
�<�ZXj�7�����[�&}��p�8�:q:���F�n�UC��?����Oݣ��hn�2�=m�8*v��O�/����������'���ۭsș�sv��ݕD�Q�qMUv��a6$���	�z��ȳ��3�Ln��cCk�,�h4�g�"����p+��Tg	hH�y�����"�����{���=�M�?{]D�!Ͷ�V IbK���Z�auwh^���S=�,��S���ZE0{l�hLX��$�g��$��*]�YB�~��l
����XH�-$#"�z���ѭ��@��@\���y�#���SFEzC�����XI?`�࠺�� ��{���ޔ䬳�#Qc׬�I�; ��-�z�ch�v:�FtVW.��7Ҥv��j*���t��2e?,t�I���Z��8$�0�o�F9��D$�]lj㭙Ӱ�L�H6����J�B\���rI�鳵N;��j�O�+�lU�5��.3)��y["@�|�䞵��V0v8$����_�����gI)�;� F����̂��\n�n��E!yĐ<��:���O��z�*��-��)��2|�,�f
b��y5������0�C?�+H��{��K��0O8.�F������|?����uX*�@�Q�[�S��I�S͐0%5&*�U�f�_Z�EY �<�!�S�X]D���K�f�����3ȧ`.|�0~�	R��_�`�_�������X)�#u(�T�r"��k<�3Li�)�]jń����U-+�2�C�����0��^d��㞅�S��3�ə��U���k{��"@I�gD�!�ȣw�������{97�b`q}�3C��t%fC��ZЁ�����c�Wf�K���D �t�����\�����7�<��"ۍ�U�
�
UP\ ؼ��E�NP�d%�;K��P�A�`��j�,�W�蟯3�jcR�I�Oت���@����)���e@�\ji�w���I��Z�+�:��Q&����jw`�)������l�����g<c�C;�{�?�����_m!p���Sn@��?��+��POqX�3|h���k�M}&��_�~s���?���M�C���7IL!z�e"��m���	�],�o���z��ټ́0�^����ƢCRm�n-�D��_�$ђ�i]b.G�F�K�$�;�r3`�����i��k2�Wo�1��ƛcA��,|��H>w�M���� h��k�$�m�k`іPꂤu�5�>������9t�C4kށ�Z�Ɵ�6y!\�7:�g�W���w��}�T�0�J^lF�@��ukj�@���m�k��7�d�:�s!E�-�y��� �X���Җ�}~������
5�ju��24��E�Y�Gy�nĞP]s���'ȣ�k�ZN���� �t�w�?YYE�.�8w�-�zs3�pc `�4)�y��cTuz��~L��|:�Ku���b��-*d��֩6�w���#==�I@���d?_ 3狝z=u�����j��@m�[��W5`,���zlFS-�ї�{�d3պ�[�W�o�oM�5��_faXU�/3QlVS,�fe�-�YO��q���M|�kW�K�:�Q�K�vf��� �	, 62���P��������N�%�´�~��pX��nĚ���&.��[���X�">i�Ƈ�x�v�����'�����E�}���#qMS��-p1W�ٞ�n"'��b�\v�b�a��������gf��qT�n�-(������d��@أ�eo]F�����3p��|x>%�U&�[~:����:�˒��Ly�� �f���g��㴌�h�x�s�	�_U��8-بU]�W�L�m���ѡsP;��˛�8��$L)�8`X,�;5Z��ܙ~/��W7]n+6�=tl��'�:c;�K1�	�/W-��\67Q�V;��Yy^��` gD��E�gd��C�؝�/7���
</a�j_���}u.W��/p�� C��l�9�?=�������ZY�MRNո�7$�X\L���OXL��v%���B��eQOۜ�� H|Zn-O��vƙ9w�|�քz+s����E���d9N�Y�A3.)���gxQ5����&� k��G����j��ȓB�⣿G��nD��s��(A�4ۄ�T�m|�����_=eWh�Z �d�����a�v��t&�B	6�;�s���A7���w�;+��o�#�L��k�:H���9���F�T�2�0-lj�aB]��9��Z�6V�*�T�M��&��,��7�����;�*�
W��/��߉��ds�O'����ί	%dU�k��df~��u�1u�!�̰R`v����X{*���I�ak��`kz��~*�8��d8d
1=s��д��=��g-�r�a��@g�5���+f�Y����7�,�+E�Ճ�����|��]�}Ab'��}\��3���m�=8@�2Å�q* ����W&�W�FI�8"Q��r/�.�a.1��V�|�25\�o�_��Q��W��'���m�6.s!���WQm��d�F_QDN#Z��0m�<R�}t彚�aÍ��O&j	�>�Mc҃�<{�(d�b";��
����.�d��2;s�-�BHjU�獴?GH�u��	/��S��GMp�imk�wlW���J���$��qQm�XM��c�!k׿�!Wfw����H�C��uiY55�&�	�g��SwD�F�·"��n�#'�����[x�|�~m0�«���S����<�|�V�h��O6�GsF�(��{N�
F�l>��g�V�{���(v/M�
V��ٽ:��i�[&߆4��D�O�t[:1v,�^�r(�
h2�Q	�t���g�n�A����6�h��_�"�
O�(���-X��F_�R&��Ȑ�����Z��~;�bj������>�Q%�3v��#�v!�c�KT����$���纩�&e��J�����fHkO�e:�L��"jE�����B��MY������>��KEFE��V�K� i��]��+�΄��'-n�����\!a�}��(x��pZ��]�S�+N�dj�
���!]SB���x; ~��E��m��-%��ִ���'�����
��"����s /��{��mǴo
b�"����0���� �=˧��v�ɒͤc�!�.�Za��8��Z)# l´�A�|Ж�'��y���81�E�śQ�E�-k�04R]��6��NsɖR���3�ga���g�!��)w�=�y*�p��iR�)z�L9��������X=�WD��8�{|B�Z����0���I�D�q�v���H��e��E��_�\m1w�kR����n�g��`��R�SF�,�O��"`�����F��f�_=�so<:"�&͊Fulg�̠�<L2����!F�����7V��;�c�xE�m�B^0#ɉ���ٞ�~O��5��f�q&��������3�rR�����v�e}��R���l�͆��X��h����|<��/֓wZ��M���P�r�+qv��F�͞�1�*'�b$-�"6P�k8o {W�S���NSn��DN`@PP��M���ȓ $�@�+%��$#B��[��H�.��%ć^Eq�C��H���(��2g���{UE�;n��2�7M,�}��܉�tf�O'���p�c���`~>�C]�&�/k��p�:���5_6#
T Z����5U���n��0��|��R
���g�+���"�
I0ɰ���.��:�j+��U��45��g�^\'�w��dbk��a�~��7�'���a��O��	� 95F����V��|����)���V�u��)��	�[_M��U��C�}(j�65'�!�!p�֬k
}�*���Y�G��z$u��ejؔ��؇!VT s% �Չ����������qar�m�[�@�yi���G]�t�Q��!rPY�D�ӫf�t�%C���ih����QF�g�H�7��*�ݔ���F|+�t�*\�, $#���m��+n��{�iþ���j̣�u���N�2#����zJ]K�{ X�#�z��F�Rp2��l�5]�Oӵ[��[y�� �C�y֫/���*���AKs�j$c��t��x;�H��B������B��^�?������/a���'��S���7��)��C* wْ����C��=���+� �����ݍ�����C���"�!>���fŢ��M�Ys�&
��y9�I��Y��EZ3��:��]o������qC�M����k��U]1y�n�!�c-�9��h��3�������z����I��_A�|��"��Z[\
Ok�S�g-!
����+�/k�"��f�D�ĩ�� Wx��K�����UU��uF�nڸ���k�r����l����_r��s�� �+�J���O8:V��'�epV����XMH�гf�����;����Pkܗ�O�������x�f�ti�~�Ǭ���9��QNl�T�d���Y7b�ͫY��T5Nw^SS90t9u�8�v%4h��4����<4��N��U���kJm�k�%*���v�+�'��o|<~��wR�5_R\�����yß�Jn��R��i%���:�ƌv@w1=�F�M�������c��@F^���q$t"v6Ek����"���SA#?��!��!x-���%`=��P|sZ��s�a8�4*��B�;z��(��4xd�'�Uj�|H�e7`��C��bVd3ʡ����Iq����aA
2���>���n�GW��߾XB�uN7���#����������$�����B�5ø9T0;��TW�F��Vx�OB�$�)n˒@����㥝�_��Rlj܄2A���
c�8��N��$���X-�ҋ'�H+��5&�IW7Ή:�����Ѻd��;m�Y�H�;���F4�r[�G��*�Z�_>O��X�9ol

����q\ k_"� V����P>���ehψ.��L�z�>䷬��(�<*�w�	���[��fw��Q
������ȟ�z�롓X��J�� (���NB� ����
���*��.�uN�i��������}��
��BU�.O@���{�/�H>c1<~���RxB���VO��`$F��p��lcѤd_��"��7�y��(���NE�J���Z�-�_SZ=�i�[�gԬ"�H�ߏ)p��NB�}a�~���{����q�X+j�v��}/��d`p�D�58�U���$�kT�({�Ů�]n�b���~3Y�0mZlA|��m��$j�!d2y��}���x����/�˿�~�ϡ�Z��x�_3��� �O�h�	���4By���z��Q�gT☌G���{{�;\�w���k�
��O��lV�XY��1�ǧ�\��tݚ�X3��WVu��j���%����m��*�� ej�^٬UV��͹".2��I�f���_hs�G�&�e�`�'�����v��{�{�z��y#1����H��$��SBm����� ��.�N���0�\Y�Y�(e����_����|8��}ۯ Q.l�}1�X�2�Euh��[R�,oХ�D�_����CϽK�� kO��C�Laٜo�}���ݒ��
O�!T�I7��J  �H�#�W0�Ɵ~j%�n��V������������K�Q��毿,���W�o^fl��_�诇��YKR��EU��M�(b��� O��H�4|R��9հ/����$�)֢�Ҵ'�8��U���4�ȊS�$}H�˰?e���c�b��d�lV*��6��A�j�촺2'v�j�/�X]��F��A�i�XѪQo��0 U�(
���rc��">J/�++��!k�@*!�"@:j��Q⚭~况�v�a��t�(�nae6�'��p�H����GNu�Ȁ:Y�'8��VK����,��3�Gk�����R�IE���"�0y�!�Δ�F��O���9�$�C����
��a��DQ�,dK������PCG2T�Zf�et�>&��RR(DH"�*AH9itǮ-M
�eA��g�|�xr�h�͇op�����0l��<=S�r_F��rV�D�ne��1u�I�坠�oQE�K<HZ���Y���\P�>~5�g����+C�*���I9�`���0K����Ƃ}���%���,ӯ���E��8*«��H+_�Kf|�7[&��?��PN��
;X/.����G>���pɿ���>��.[�|����z�7�]?*K�1���JI��_v׫��k�*���%�?˂�ko|�y/�������>���j<,G�������Ύ��b���Ϸ��x=N�d9��P"3Q�}��˯��k[u�����1rRcv��X��;�\, ��bF���(݆t6��)�UFl��E�RBW+�Q�b � ����}4F��/g�5&a1�Iu>���Y���ac�q`ڊ<��
	��[���.Z5K-D98�
��ůeE�����b���˧&�&�ZV��XS}w��Bs|�P����%���,�a�qQ3�n]�.v��5�) ��e�C)}���]|=����Y�4�R��?|rx(�8��s�Y&�Ө��މ�pu��+�������B�E{X�@c)j�-rg�A���� oAs�c�]����R�y���e�P��.��͑��C�(��9w�L�4���&;�OD��QRnH�>�C��A?��2'C���1h�Q�_	�A��.��{�^�r���<�Od�y��r6�����O�b�|T��b�oX���-�c���v
��E���'W�$������t�n��[�Ū���������'E�*X�W!��!��� ��=���;�fNv�{���j�\\Z�a!�r�ŻP�PV��ل��;�!�h1{��)�7�� ��D���'�t{�ږ3�I�����X�K���+���M�=��0�3���e&x�@�^�0�9����8��6�	*uЁ�� P���VFU!�_~"B�T�����6��Q�<a�q�\z�+�������/1%�2����)I�Ί+�(�I-Hb���;�t�Q���u�	��D���K�i�����P�X�h	���w�j���JyKrDļݶ}��1�b{�D{E��pbFz�׏}jwp[ز��2PP��8�p�*��*��`)Z�Kwș�#,�2+p��l3�;'j�n/Y*OXLEw���C�7I���2� r������o���cZP���0�^�M�"&Ť6>cڢ���G�g>��n��Ak��rq�����s�M�, w)�C�ZGM��
Y�U�}���u ��ʬ���@5_`c������v��]p��ӻ<vH�4��l�%����5N�afw��]��m�����з���n,��?���7h�����K �|a[�ޛX�&���A�иÇ@KS��l�F��h�5�3
9m�(�Ã�C��^5�cƞs��Q��a�)x�ŭB�	���4��hw�ǘ[�.?K�� û�wNQ5���b�٠o�"sPE�: ���m[	��d�J�,2�&��
��'�8	
�}0f8�1�U9/I���d�j��6�u��Ĺv��*4���Q�n�w����@t�\�ljO��٤J����D�8)4�:���L��V��Ad���V���Hją�a�!�rl��r�? ����x=�<��'d\�ޙ�3�+���*���R���ԅ�M�pU�
IE@�"�9@\wV�׊�⢕B3���@�^�����	B��q<�"ltb�����p�����qV �N5z��4����1�܍,���/�  ?(Vۭ{Yh����z�Tc$b3P_�
fIw܄x<��:`��>"%�ȷ���}IЀܕ���"��	B ���V��O�����'��{ȶ
�ř_L�#�!ղ��f{��"��0锺�wr�'U���VԔ]&M���^cH3����~6�r�*!_�BI�����l���'+ݰ�?��Y.�Rѧ\������ba����f��)���_�Z��?�6I�wK�D2���v7`�4,9>�"*^��]�Y|�?33VH���_�LY]3 |�㆐��n�����Z6�㌰��Dc�t���`CW�����z�3塴�I����R��Y�,����߆A33)_���������Uz�}���l�G���J<�ʎ�y�ݵ����R�TT��{��Ll]%�G.
TM��0x��]�x5liB9D�tT�=��@g�,`��l�~�/�� e�֑
�u]]ֲ��~�]���9*����!D��p`׃G	ߑG>�R��c��y3�x����-�h$�@������M���4��jv��p��=&p7� �b��w1�ɱ����ܝp����{j�u{2�H+�	xeӆ���͉#�^����"����m9љ��B�i�L��������jW �Q���W�3�H$�3���)������c@^�~��A��ע��Vo�!Ñ������Hخ=�pt������
��V ˪�:#A7&�h3��>�/B�޳g�܃�����K����P���?SM�Wta)��|!3��0n��Ըe��o��n��W��f�����k0S��y�����٤�Hju*���a��͝����ӥS'cf�q��@b�SO����郵7)ē��N�i�1���w�ӌ���wd-��Z��Cv�`�o��^�9Z��U�7b/1��x��Yo�I����s����ad�O��8�=�B���Vp�;�pfW�陥���X- q���l� ���0W���>�P��2���;)����_�V�	+]�$���zopd@�����9#��7Ж�O'�D�/g�aCu>�����K��H�U϶[�����z���q�wmC�����d|}p�#��ʝk�I=Iso��3W���a ?�B�'�ܔ�����)Mr��0�RZ ׁ����2].�O������*�`�1%�ebˆ��Ӌ�E�
�E�S*N��B�IkS���s�Bc
�}��LxT���]v�a�[@�I��CO� (?��7���T
���/St�@"�<-�s<E��ؿ|���)���%��[IYi�q�k8oU�K$A�I` Fd�����{�JX3� }���r8b��������jE!؂-݉]!vHV����+��Bn�a����0f�-�	x c'k�{Cj�����2j����]4�h��]�2��ӦZ~n�t�W#�� �����w����������;�ZY���b����F/��B�Z�7y�M�m˸�4ː�h1�z����;��µ����ZP�)_;B����zn��{Ǫ��upq��cҺl���t�-�n�3��������������En���v�`%y;����kߵ�_�u���E�s�������Y��R5��2jY�R�IIh��π??|��\��B,-k�x?fQ��W�Y�az)m��ajy5Q�IO�KOy/$�ƾ���
�jdC\YE^m<�i�JVA5p�U�^�&��Ϊ=(nM�iʎ�*ű�'ͩ���ꍉ��!ޅz��6h�;Ԧ���D;3��H({}aj���FG<FD�5��Z�}D	��[jm��v���`�v T���`��͌�f���j&��q�lt�!&��4�����Rڴ�0/�x~��b�5$>���2��ƙ吥��yv�Qxfo畈sj:�x��݂�N]_n�t�3J���"�c�f����f�9�g>�@���cC���q�W���������ɻE��h�,6�{I)K�!�/�b~}���� W�y��kd	���k�`����60�I��/:�Ʈ�*maa>ϋѯ=C�/~�2�_R�M�Y����y����!�L}����ܞC�=�<��#
G
5���ަ���_x
��V�������b�&"�oSک�{�h�la���B�փ�x`�q|��D��V-�h����O�C��V܃��N$��u�Q)�����}<h'���J?��+]�OV<#�p�S����Q��H���dS��ws¢<���-��Ƭesu��@���L@w�p�블S����4�!f��E[�$���ō�AoO��8N�8T��\;�Ϥ�?;�u>C��(=��I���ܮ���[!q���}J��0�Qŷm����]��
��������NO�x ɄC���{P�r�敗Alϴ��
���([���%����#q���&����W��T bE:&�m���is�5�� � d=bf��$k�0hY����SJ3.�'nd�E ��y�W_mHB�2������c~ G�H�)
r�&��|���kNX<L��9�&(-K�N8n%eL;��Cj��Ѻ2�B5��U%?<[�$R�X���(��^�p����%����k��k��+-=��<]��ͲB�,��.��un���)	==^[6�V����v�f��+sUٓ )B��)��-"F�Z��:��k|���)6���ˬ01�|��8謖��ɮ�#��4�;��˸B)�dq�R�T}3�������ب�/�����uCU��<�-�B��=�����y���Y��y����~����Dܪ���p�<�h3�C�,
�r�Ǿ���*W�(;�=�I���l!R���T���% �v���G ���'@��Y�(�oQ`j���Y;d�ZR�w�u9�4u��*�:|@.
���#�#4�,*Q;/��t\1���Oؕ���11<O.��1���uw�e�}_���,�jɪ��Pv½4 �b��ɚZi���*��,|���2�D���_��
]�̾��=�KD��kb���᙭g��^ܙ�?�b�?�(����F���g�#h�`C�W�=�6�u]��Ry0����Zv�quG�NC�n���=\.z{���ߎ�-��x	Li��UU�/D�ls&�C^&��D�Q�c�}�ηJu�5ᩭN*#|?��'Lr�8W����		٭-J��AZ�{�����V�U�VH�J�G�/�G#g������3uدa�p��{��uO�>t�b�Lч���3{�"O6��t,Y'*��	��Y�dp̭Z�`��>�
�F�f/h-�9)'���n�������%��|�Վ����~�>��Z��z�J
f8݀�u�~��6�[	���xE�g��.w#��
K����+�s���5�7h,��O��MN��b��:�'�e����!(5�ϩ3ξ+�2�����7���G�4Hrg�g�K�j�D7�!�aץ3i�'�T<uqo�xM	2�N��R3�|�:��X��r�V1o�w��Y3�[۝a�6�'a��٠����,}b�%Df�]
pϦ	��y_12г���Qrfi�7&���K[��ԪrvJ	���ж-���j���!��l�w�u�2kU�ʖlX?)��s]�
&{1���a1!t[�rZ�bL'����ۺ���V�`lm] 1J�!Xa1��}�5�B���#Q�V�"pmL-��7A�2��r��mqu����T��1��6mpM��$� vI����ǂ�b�O��+
�gL
�񦪣� c���r=���X�!èf�[w���k/� RjLo߿�ʃH�k�'*��=����Y_&[��	G�(8>	��#.��q���u���>���
G�"�����XwE���`	�h��#/^�K�_J��%.���jx���C�F�+ӟӡ!�����RG�����f���9��
�0V�Ȣ��wWR����Bo����ܸ�\��5�I����%�Y�����ӨUP�͆��jR��@�)�lQ8-�|���\��s���L������݂���*�b¦��n9_��P�鵍��va�/�,9wF�:��>�Ї�mqa�$x�RZ���]�+K�@�|&BN�6�n?�&�w*��r�40�=�Q}b>��X0C�n�Ю�
��{.[�)L�m��Ԟ�|��+<�3Zu�Pפt9�6� 5u'\��0��{�Z����d�ʓ�"|w�,%�*����h�1��R�'m��mۏ���k$�ݏY�w�K	>��:�=�gk�3�k���0؇��:ޜa3
�*5�Zj�r��d�%�b��0�R�a+�<���S
�� �e������vJ5��B�w��ͦ�[�Mg+��D{�Y���+������y5J��d�9���?�d>Z!Ev�fgz�������CIKF?��3�K8IJ���͚(o#q-zD�z륤��*���{�ڭ��B�m&�"����]��k�T�������N�9z�t�%Β^�cA:��?%�H6�Vi�a��-+��.�T��K��f���?�dK����+j�[�U���J��W�cf0c)��;����P$��Y�n� g��!��!o[T-�	���Wr��+�`�B�4��US�^���]���P[Q��Ҭp���}��:d��}��
�w�W��b'�r��~�.P���jZ������X�rl�p���AhO8�b���lܤ��j4sVX*�i��*U%a���8�j���Q^��6�֬�2
���x�YN5+޿�R�T��K� ��(k�������*&����l̤�%�K@;L�A��p�b���|�]��֟t!���\-*2r�?3����&�
Y��%�� �������6U�O��\�U��b#�'�O���\���^�	%x=�I�_��9-+7<~�!�-1Mx[�X���BJ�6AE�]�U�.k�̾��#���XA��;^m2�4/�HSh.Ę��x�e"�C¹
��J̸Q<����2�ғY�RLH+�5�A�L=�$m֝z<Z�ȥ������u^.�XUy0������y�����,Ψ}'�������%|}��	ًh���$1�����^<@�hHt줾,Ȯ��W�|B,a�	��
��V�J���ʐ7w'���dV'��`�>z�.���vq��*�����&d������w!a2NQ����B��<�\+�ʐ9��~����\�d��5��qѰ.�O{�恲6�q��lJ��C�T\����~k�/�P���ן��噘>9`�5&n'*ө�	(C��Q\� T�'��F$,
���Z���@��?���������� ������5�=�c������V�l��A��v�	`7���/2o�;C(����8��r��n��yh��f��[W�#�BM �9M-£�٨~Xį�>�P�@_����gTn�si� v&\V�"'N��D�u��[����r���P0�����wq�q��$'I5�7�,!�dBP)_1���G?�)T��2j�k>��eG��}�c����f���h����a�ڝ�u�{7��NR���L�!k[vՍ�S��2T5��T��L^��gە��)�A#u��nY�6��q|y���%��W w��WqH*%*����o��r��䙃�q9
3�b�ҭ����*���� "Y�ա��ęf����U\�����&0*�Mrܙ0o�؀�~"�I%��b�}n6;����`�Ax�M�vv ������b�?U��o�������=1�WG~��c�"�3�d�����]���b-����O�iiڄn��Hz�/c�e�{	�uc��N�ۈ�Y�ls;��E��0X����2��q�5� ׶?<�U,�/RV��l�@�(͈+��ڮ���@���6�V6K*�Jܝ���L�����WҌpئ� ��#����e@pQ$$��b�д������i|����R��)L�����x޿�+�M��WG폧,1#x9&l38��:��S�'B�<�s*�-�������+� �Q纝���P�+-k�B�.�moni����#�=Od�*�p4 �<t�
DMP3��M=�w%^$�r�q<.�n<�����XMO;�����|]&;��Y�K{P��1��HvT`�B}Z���ys����[T�.�����YW�7�b��*5�I2��;���Rn�b�s _���gv	������fl:|A�gG�����O\Kz��w�P?�0���x)g�23�6�z
���Ǒ�ҏ��#���&�(cl�I�St�B�< k�AZ ��h5��?IX�$�_�"Gx�����ؒ*�"h��^?z\�R���%<�#�t�J����<� |('(�O��S4�hU�{ Fm�A.#��@��;vTz�?��X��XF����H��}���E�t�k��r�@������� o�m��;���;�p��25����D�����Q��+��7�p�%���#-���T�t�	�_#j!�=I�_c�[!���U�P���
�ֲ��7f.��rbs��-U�* ����N��6/�_�zC�`��\T0�':ߡ�����'�u�'�h�� ́v�@oߒ�Щ�P]�G�MM11�wR�5C��^z�8�������V_Qh�[8��Q6w;��\-�󴓳R�6����%�����|oV��g�.�w�*��M���AE�e���T ;�>����z��}�M�ADN��T��u�J<N~CZJ�址?#	D�d�ܑ�,!Ru%+Wz@(d��3�OB�裢:Kxg@݄�&����$%Vt�� �/��PT�ԭYD�-bqB�rH-��.01����{�Ww[��x$�LW�q�<sb)E�$��Yj��$����B �Q�.�θ�<�uޡ��t������L[��>l�0i���7��qY�s0?.\]�gء:���7ޜ�F�*;M���ҷ�ƌ�T���2��4���5	G��k��$S��\���� bKy,�;@�P2Ͷ__5�����AAӭmQ$�6�qr�"���a&�'��^'��x?\�z˥0qIMz�XN�Krm<�N�&ϟ�L�Ӈ2=�`)��U�U�\�M�;��\��ql���n���&x�U<m4΁��j���	]&�t�AW���W&-��P�Y1:�7"�~p^��#��|ө,i���dp<��4��BR�"��ɤ�<AN�/�銳�2f[�_�=���=F5�c�B�ٛ�%O�bv��u���4B��FǶ��.�7��n+�h5�Z�hH�*s�0W[�$�4"��2�>�l�P���
�j�'�T�j�!�x�N�0hҧ�s~?T Z�]:bhCG�zg�C�s("\���K@�D_��K��W��b]E-����<�����x��s�>a��_(0�'[&u���%oU����|������CYW���l@��ۖ+H��,R�����q��9�/�,��;e�W~HU��|��n��7�?{�)bq�ܖ��
�wsw�D�T��Z��C�&���+S�I=��v�^"��Z���Wr�MD��$SZ�����.
�h[�7�r�M]�6��e�O�0V��Ӷ8ϕ�J����̔�B�3~��7�aEiA�kc�a���Y��r�zN��Jx.e��s�(�]�����JZO�S�g��O�Z�.Ttp���U��ǃ�+���BX��z +6�iA�����m	Nj�
��z�)/�f+EѢ@���ڬ	A����d]x��Nwu�(u\��%<4�J���*��Ӂ	�<�<jr�NgD�d��=0�D��(�$3T[�10q� ґ���s2�E�y�C��r�,Z�h87J3q�è*��=�����Z�g� P	�W�[�b�o�1~Ȝ��~��9Z��8�k�h#^�Ć[�5��`<U���J�6s�2i�
lѰ�t�йd�w|��L)���+4mx�l����@w��)E] ���2������Y��hho[oL���M[�[�p�_�2.0���Z*�f���7�
�������ω:+A��?I�.��v�Lqn=�ָ�E��B��j�A�̓�K��"��$z�?c$�h��'�wˀ�ݽ�E~�V�]9��9pW��[���T���с2�r:-���eb�R%]B��ќ�L�}�u�-��wb����=q��3�˷IE֏��1��/�:O.ʳ,�Db��D�JV��om��8���;֍Z��柉Lөz�4w[`($Ѱ�j�r���:E&��'�F!�[#���b�.dI�Va������q���E�N�]�fQ�J��3q���紜�>͗�X�0?����$�z�u��_6�1,��e�cV�#nPEz���n�f�pg�IHc0J�R�"�Ԩ�b��[�+�eU������>XP��J����g��������.q랶	���3bc�qc	�Ʌ��Æ� ��8{L� (��Y�c-���k�ħ��;�=��Ie�`��3�@)WЂ��d5�]	�@�Y��L��5G������|��
�#�rڄ��r�F���>=��2	�,�ʹ �QM{,nX韏٘�aR�76A�PfFaB�Ŝ�G�ּ`	58pr�ޓ���7�z�515+)�t�>�K����S��O��£�ң���
g�0(%���� ��gr\���#g#�xzn�Z"k��l�Խ�_a��A�Td�@���RXHQ��B8��S�~�p	��%G0���{��J^�>����v���B֬v���9�38�" Zv����?z���K��<O�V$*��i���光��i$K�e�Ɩ�1l��Z��D����L��i�s���d�aS���N���^�z���T��W1�i����L�pF�|��%�O���+�Ƀ=*�&��� ����%�iw?�8��*�~zonw}�(�"���0��z�Ysz��Tܢ���l|��x��QŐ�����ا�]a�
p��z�Ǽ�0�Cs�J�L�V�5�-���km#�k�%�T�@�0���U��<�Br�d�����	�1��^�[��3������M4m�b|� �:��*+�K�%���r�_� O[Vn�
l~�ּ��e����q�j���8H$,�Gҩ~��wJY>�O
�j*��0�7W�#���ed�߸ZhȮ�+� �I]
ǩI.�� ӣ���2��6���%l���o'!t��}�-ޚ�wRT񛝺�"D9�	����]�7�O
�}�8�" �"񌡷R�v�9D��}��KGj�X?8��A��oU����,�m�����ѻ�֝��yR���$%��Lh���s�ͤ�^zfV�6]�����ʹ���l#�=�`f �#[��ß%	o���J��n\�5��PR1���H�B(@�(� ��h~0##��{��jL��G�#$=)�]����7�ܑX��a����|`��d�S�0���w��cd�Ql�F�B`L	�"��&�j�e�����.İ�N+# S5r��6��R>*fU�Q+jS�I���TN�(0ۼ�m���U��5�_�6��Ծ��῾)4 \��k�1���5h��b#���F̀��^g��&���C�E�%δr�4L�j������E��A|0e��2�\
.���Jy͛D�2f
��n��!b�ơ���\\���_�e�wa��MB��D��� _���ڈnJ֕�ͻ/���{��(�*�Z�,7����C�I�NQ�ν�fx� ��ƐA�=1�z��4~���:�<-Mt���&���:�9�'Z��|�
���4��/����{R^� �a��G6����ƳSV�f�,���utp3�|��N�:Y�HExZHU��[�q�BBr��sVCތ�Xy�_�U�2;	аu�$���>G���b��ɽ�7�Y��IƼ��B�i�-l)�Mlz).s<I]�տ�̀����빼�Q��x�����q�N&U�Pȍ�r!�i�N'R@+�Yr�2���3��/ʻf���m�&f�c�w�r+�~?�V窯�b޻����ҹ�CKM$1�o�\���a��v��W[����핝�xB� f�&����~V��~9��=�s������ػ���8"�	)e�]��m� s���T��8�����wY�)�9'��2]�{�Ё��+��-��%DE���k��F��0wi��ޘ��v�Z��Y|2����tYY�z��gXֈ^����mѯ�d$C$�x3�5A��%+F����5�Xg��^h�i�J��[���<6��`��)|������Yd>�.NNs��8����= �P}�����f�Z�I����αQ7y~nr���v�,ȭ9bb��!{�N�{^��ר�O�6g��%�"Wiz��7.�
]��{�m�N�*�#*�{]��_�Uiu�`��47��Iɱ=Jmwmw�l&_�x郇dQ�K�wծ��a'[�;���*�wqȫK���}�G\�W�;�nVc�X�
p�[5�	HL�B
x��~+���k�p"P�=�Z�g�>�[��퀧�>1�1|`�'��fUha5����مV��W&9��/FM!�nHu�
�=F��"x$�
"���o�����Tq���5֋��X���0�����g�����FA�a7��э�8��W�j��W ����9�QU�(�3�szXv�Up3�y��tq��U~kE��+����dj��,�b��2�	y8��7y
'���L��2ηڤDhL�O�,Q6H|ҁ����0r��l�4:ijl$���x̀��q��� �4���^K껗nx	�6pX� �2*�='��>U�A��?��� cZ���	{��t��Zr
�hc<��ALs�t�w���K��h��z��P���2}����0Z� �`��TAq�P���gnx$]Ao���;�$\ԢX��cڠ=٣�.��~>\�bԌ��6M�����:�'�2X)b2ǘ�=�Gm���/���ɿ�ڜ�Sit�bD��B2c7��YX�����)�@c0�ԅ^�:�F>��T���&?yf�ܱ͊j�z��-N"WJP{ͤ�; �䤒�n#��Մ�����+lH�RhQ��$�~/^�����T��|��_�DW�>:�����3�>K���S´j��s�8X+?��T� c���1Ea�O ���M�7'���h�X�'q�K��m�#��=f�3�2SRo����̦RY��9o�!I�}b3KS蕡���]���3dED9K406@�$o���j߭��"�3�������/g~4x��`�֏�b(�\1́3�5Z��l�kL��<�E�V��p� [� ��s7nGⱪb�\�3OB��鯈� ��d������gJ�[ ��JFp���9=�b��P�I�؂�g�2)q�ꑗ����w4�<'sw$����ߔ	(k !-�Q�1�R��>�A�e���p�5���ja<%;B�L2�q���C���[�A$��Jƅ�ŗ�MҒL<�(nJ�C���+JJ.,� ��qF�3�5g�;.iHa������n��Hz�+!�_J> w��������-��lC(o�j
�|�E�ٛ�bYO=��
+������ʞKn�����%�ȲM����6��zz�4t�?!�fH�"H9[��#�;��{F��i���=g4���?��,����|B�_��͎�-�`O�ϫ��bif&�O�B��8�՚g�լ3-E��+� ��n���^}���2e���`O�jl��/���¿�0G�V.�4"��ڒ�uf3$V�ޯׁ�.���y�}�Y>�A��j� M�>ڡ3�#a/�޿߉>��7�N�6e�ӂ���M�eq*il���R�8s������@���^��>:g)���i�#B�֢M��IOc�_E|B�{�@д������ݫ��O��f�S8��c"�aFy������FX�N���\G��i���֨x���l"SHo )��x�ت�������1�C�#cHS�ט{nc�`�χ�-��Q|�׶�Uߞ_t�^8�W�8
��	�'�V���+�ɚL�YX8�\�Z%)@�c3����ɦ/�l� �҃'�i�g�݈���^(������{C�0�FٯH}�#�_����Ϻ!^yP����X+j�)��3:yn�\���X$D\���	�"G�n�	w�+��Mk;\7�����[��.2!��>4�����̜�3g��76uV��V[��#��(����q��ŨuksNJmcz����N|��6�,E[֣9�a�7�C���G�l�J�&	�D������P8���t#�W�"V��3g��7O����@�(����;����v�⺟l�"���Z'3����(f��uP�J�A�ZU�d#����7��t��69�u�pFm{��f�6�������9m��f��)���_#�NOI�˵?f���
��4�B{��������&�Q�e ��� �y�~y���FH�(��d�-����
��[Y�uչ�_��:��p�$A�8�K�*L�5�p�._:�}�{>[��&�p�I	Kf,����-����am���U��R�Qҽ�=������}W�;�#�
1�fK��F���H��gƿ�}���2A{���؉?��{�:��qY)�(�+h�ē0(|U� '��ͷ+��5lE���rBU��f[ �~�� �Xͫ71�.�~>XF=��e��zk\�l١v�T1$��%bI��ӽ�a��w!�BJ �e���������Ѭn&5�����|8���X�	~$��yxݽ�?�BGbҋ�s�@���V��p�f��;����"���Q��Uq �j�"���Վ��6l����g9�c0������O�O|6ث��	K���RN�?�A�{Q������&έ_0c4����F������.'��i����/��<>V:��ހu��و�&e��L҂�J����ܘ!,���+����v�u*0yol�����X��Y��է��ea�L��0�Q��V�u%E�Ht�~kLv�.r�,\yk)׊�4ON�1|��q��(r~�xc��×���{1 .E݃�e�j�<"3m�߭3� ���ߧ�i@�7*.C3�֚ZPո�A�7�dռ[�5��E]s<Ss!QG� "%P�g{�.���^�E�1�+˺�q
bg_U�#�e�m8���>�g�D�2�%�����~�i�z�ʶDŁG5uE�e���`	�\���Z&�3�92���������Jlں������ռT�,�l��}�W��j��w���6���7��[%:�=r5��vU�
]]�f��LN��XՎ��0�*Tg�k���[O��0B�\̳Ƈ)���E�������ą$���Ajc3
r�^>��wL����je[��;��ٚ_n���u.�&a��)শ�H3l�,8��O�I�A���L���|ȓ��C}��Ҷ>�SG��R���:c�e�f�n��L#���{���]�μg�*��]�K�o秈���]��CV�mEQ?�4��r��"��c(@3���[`�4[�sr}�o�t#9S�+��Q�?>����)kw��;*S(��>�flN��bFfp�w��'_.܏[�<�g��(2k�=no����Tv�l���%oT���K렇�� �a�ӣ�$�Bvɚ@�e'�yH���|�p-���^9Q2{�������L�K�j��JuB���1ƕ�!�N��-m�	u{�)1��Tf�|%8�m`W~�\J]DM��e++AK&ئ��5g���D�*I��pHʷ�������F!��v��)���4Q��c!����p����m�
��w�Vޫ&5I���1�-��+"����\�,Yn�0���*п鯐b��U�Ƌ�Q�Z'� ���eJl�z{�Y�2v����԰%J�g�bIg��͈��^�ɯ�	AB�YΛ�ͣ��4׫7P�����j�����H���
5�6�¨�����0�o���~5;�=��Zh-�ͬ����^�u��!��H��Ø����/��j�s�Bf���CF�!{c�G��.k�sSBl��:7�
��ޜ��a�Uj��w=�f(��8���|9J]�������r.��h�L���G�888d�	�F02R�LyN����u����>{����jp�I����+���N�x���Vyi��Lh�჌H0���%����:�Yd�I��j����D����,"���a�4g�$W�]n���t;���d���C-���K^=66^ѿ��M$+���=mza��;�"�_��Q:��4�C�N�2S_�+c��9��z�P����=fP�>
��)�e-hk+u�6՞.R����{���ƻ�(r�{�ce��D�BdD��U?�\o��Z:a�!�R���[���6��Q�R��;�������tEz��_1��R �}�ﾣ�^�P��I�u��G�Y�p[P�Xsy:iJXA(���G��ozk��R�τ,.⭫�k�����$����4�VΨ�F�ҾP�i*v�J��_7xd�fJV��aE[�^O:��(W+(&Z�*Ux^��Y�Ka��ڪK��qr��Ͻ"RK�0m��Vm��x�2��*��F-Y�8Y��{-opE��_˰^}�~
�Ы�)���08�y3������"=Ϛyx��2�܎������b͒�d����^0�KCS�ɇ�r�+�:g�����H�����g����#�����£H �HP�=�@��c �% �o:5�*�8��;� �]�{�CțB� =��C�1+�u|ڑ�����f�p ?s�`��jQn��w�d ��+ΦVU�%��w��4n����V��!G��x�;���gf�!4�?ȯ�GX'ϯё���3�9��P���ޘ`��!*i&ńs4�[��h�Ńv�����YY�N�evP�S��������Zq������4���:��iS�'�~�σ��ۧ#p�aa����p����	I7§�A.C�Q�DkRi
���XU��x��˿����+�#�����=�E�Տ�QJ'�#">�K���p�1�a���]{P�v�_g��	�ŵպ�c-a��}��5E;�A�PQ�O� &o �k<���Ի�������t�`�
I�K�i��ɪIVi�̪P�O�x�D��\�c� ��fXx�QbG��<�d�$�u�0������<i�:���E�P{�H� TL�"�ߕ�ޒ�p�׆��+����@ �!ZU�b�p���ޛ��8�����G��]��қ�Ld3~�}_vz	�?�h kQ����Q�47������Z��e�]ƈ����8JϒIT��"U�>]]_yŲt�M�+��2jM��n�}^
�d,	�U���r���η8y��Ivm�k��C
�(������KQ=�7Bu���>�6踿��o�"��?}e�0,��]���b��1����N�g��\��z���G��q��;>ݕbW�� �3��(<�5��n��M~_�y�a��J�����յP�����4�crdu�5��c��A$��,�����齶�\|W#̐��U�r�@h�y�o�U{;Vĥ��O��U"����PX���WʤQ�����w�?������Y�tx��K�rj��X}��8�~�C�Qq˧qR���D�)���[i�+�@�>�&վ��t�zY��IIZ7�OK�f��רF?#�pA�P�E��S'��i`~����n{�q��K����.�?��z�������w)�RbZ�h�2G%� e!zB���"9����Kt6ok��E�(��`^��1?FK�F����Si$A1�1?�^��j>�<3H;�yH��N��
����f)��Fs)@G�rه�Jq!͎���
�*c`�~�W�~�cܗQ�׍.SD�5Ӫ�����H�T����^��=��p̸�(���=�D�g]B����:���]��˔�k�������V:^te���> ��"y�{�/FQ����޷%���^S�(�O�x�q�(��͑cw�5#k��	�ƴNq���í ^�$���vö�E^ka��oW�.���ڏ��/���#���z�w�BmCf�7tFkq
�ޏ�Q�y�鄥ۀ�-6�-��T�.�O� ʂ���8�;�w�ԉB!����K�敺r[T��a6ˤ�Kg�u���%8輆�G1�����g������q�H�������4�6��Pp�/�7ai'{69u���&�H{?on�@����#>�*d."j���� #�,,;}#F����9�ãx�^����4RW끽���bO��|pE�7����R���c���bҺ��J���V�n0'��ho/R%xI�T#'����_Ei]I��f�y�����*�3�'ˊ�5�Vs �G2�cV��iI�Ѭ�G	�'Ƞt�l�p%��/*!��lx~"���׊�-���T"ͽ��'��+1���b��r�e�{�[�&A�)#>��l/³Cڅ��D��>���ݜ�3Aca#x
wӻ8�x])��������߃�ȣ���x`N��ҤC��T���gT5��b��$>��{��nۿi}�,���`���xl�K�s�.�ޭ�k����	�KR�,J.cP�� ��l%�'X!l)�a�t�~ @��զ
�)Qi�O�p 䌣�R6� �˿����V��?��t�2���y�����EX�;pE�vAk̟�|Q��ȼ�/��]RΜ:�Ul��l�1s@k��%��N��JI*JxyҺۀ�C%������m�˻��wH	|�_3��D�`u� ?@E�<y�����6M����fd,��w.d.؄���ת@ȭ�)Fh�@�Z�DX|1$?��^�@O�F�ƌ}S2��Je]#hI��ÊD#o��?�L����߮�;���=Q�"���$��f�bZ�����.�=!���PD5��<�V�/�|8��8�H�:��x;�7��s��c-�ܧ����BD�c�^�q{�R�Ӫ�m2�S��gaC'�-&��*q�����#	Bj�����WZL$�3��n���yI4��	i \��e)������l��`s�F?���n�ƃS2���u��_�L�Ή4�a�Z�&�C`���H��$�%�gG�R��Zf��.���ɞHf:�ۢ���������Kg�X=�V�+^d�^X��g;ِ�?��`	�А��,���&�~i*�r~QD+\=V��C,��G�6��w �Zh�n"��������Є��A��~{���9��/��|�]�~B2�wv����vd*Ъ�e���:1_"��k�����r�3�J�J-�WB��/�V�˧K�ȡh���[���fz���OH�[k�=�{�(��{�nZ�Rأ$�|A�b�����꫊ֹn���RdB���j;p4e.���W`��b��m�|=������n<$����<�1R�E�S������^����F'�g��!�_��<�J/�(�P�0G��d%�6bb�E*p��Uz�փΆ�a������ة��ys$6��ۄ#>]>\ �s� R�P�+��֟��o5Tc���k���A_�$�f�ˡ[|BU��h��#kBՆ-M�$r�˃P�Z�1S�qưIAi�.�@�N�=J��0�Vw]a�YWj�k��;fh��
�'���ыU�f���d�evڗO:5D��7�-~�������$-�E�|I�����߭�0R����I��*�F9�z�-s*f�\�Ew���d+���c�RL��$��39�5@�Mo5I���ҽ�J���V����vM#���hYl� �ݜ�wI��Ƞ�(�/�d^�e�{���O�.'h�8��-����SJ�G;3�)Yt1E!E�q!ש��M����j%A5��L,�ǯD����ˇ���2���5��D����A�7�$�+�Û6��Q:�� h�6^��n����g0LЗ*�vI\������#E��̈́�!#g�8�"h��������rŇzS�c��$1ߠ��֜)��{����������
'�y��M�!�:�g��x�F�f����i�9���%C���kh�:�r���#��3�E�8�p �5��`2W��|���t��R�8��A���'
˫�'u�����/a����-�y>�lJ71��&@�X}m�{ȫ��r�:#i��zU�gV�PSs�ͦ�<�"ǳ08�����Eb��M��C��,stGgM&Dg��U��%J(��:,@�v~�m"����'��l2E�S�% G.�������(�|��@~�?b�ɜ���9� �y��0�;2�x+���"��<�2�<K�?��՝�V��2ׁT�bE�P椽Z���M��5'|�����->|n�zrᇫ�-�^`W��Lk����ȃ�q��S�;p2M������<ts��L)�2s�6����r(�
�o8-���V���hW�Ȅ9FxB����[�XJ��֐�8��j��*�,�~��4�Ow�����B`j�c��BVc4�|�[B;��Kc�c��U��Ǡ��]�[U�p�������}٦�J������/{�	�r�*���V[/g�Ѯ,�����vOL@��!��B��_
�z�f�!9�MJ��UvL(1		.,�|	�Od��=#�*�?w��\D�?���b�>�7��M�G&��GH�5L�X-VBd~��QشO� "��_s�'ԙ���mBp�㵑��4���@�ڞ�ʪ�'�pN�E_��W�gR�_�X�o���K��/>$z�m���;��%m�W��[�A/��C���.��oH3p/p�y	���W�6c�"����ĵ1:�Y�b>����vHq��Q�-ᡟ3���L�����v]�b��H�/+o���O
�����d�qg���Q=��8c� ���2�ػX�F�dmߜY܏F�Oa-���/���_���` �T	V�)xN0TF��_�B���z&h�Q�2��[ȗ#�[���ܕ�8��T�c��~��w8���cソj?ޢ�r��ַ�b�_�'�H���zh׶[l3�|�$䨘�t�@�3 ��2K	//�����D!��>Gܽ%Ȉס�O��9APPoCh�
��c��'cS���_-�jR�9������7�]7�Y���ň���\�M\X4L+�i_���tq9���ڂz��\`�Yj�Z�	u��!p0���ډ���.[8'H'yVǄ9`��ç��%�9dS��)��u���#�m�W
F��y�$�/�E���l`PE��(�8��@²��%y7m�Cb���_�g>���q��/��¢��7��ma)�G����b�D�J�?�S��3��Q��K�l|_5m�\aaǘ�Q_���'�Os֛�v<�}8���� �$�\�/�6�Se4`�B�]|^�A�np�q�f��%�1�lS�C�ت�MvpL�������ؽL��}�Y���t���7�=�*7�k���w���x�K�3T�Y���������)�K����'ಢ�SV��Eg��!�}­u��7!Vԗ7��\wye"��'}��?@@��V�=���%l�i�g�C�Ƀ���~��Ě8˥(�,����x��?�F�}�[�vk�ډ<������	������.6z�1k[�W��oMNt/�e'��i�`k�6�|}$��زf	a
t�A^�| (��LjF�!�}w���h,
�@�II������v�w����>����Ti�.ؼ���Ϭy��d�A�Ow�;�>�!����8�rn��+Uz��K�({X�.ę�W�j��Rc07�Qt�ؘ�uP�m�r'Y�#��nI�����F���&q�Ya��ޟ0`m�@��G�^[�P:Mw3
tA ���o�2n�G{�z*��y��Ɗora��:;8AN��ڀ��u��ut���s���qz��Uˁ��{o�d�r[��oI�YW�%�P�=	#���{@Y�*C���a/ %������+3���Ra�B!��8��L�'W	��?����=��C(A#��ڴn�`��a�AQ�v��7Zx�aȜ�/���x�ןr��b�R\gA�m3i ���?ZJy�Q�I|P �!�WZ�^w��T���o�ڥȼhI�#s亿�0�5஬�EZI�wx�.W�M=O��t�7�*��UFlN��Ỽ*t��؈���/-?n�n͇QЕ����[���c,/�Nf����J�LR��D�P+��_6V2�Dz@�����[��\�g�����8��KEA�%k� ��6�����*�4P��������c��um1��ؖ�Dt6S�.�L��wF��M�1ߊp�!�uV/;HU:����6𱪛�sl���i@�ն[u�F��V�0����膟��9!�	Qn��2�n��U)�����]bh���S.����K���Y/�L7�K't��Jyo�?�<A���f��f���F�,U��b�kԅo��v�T�$�i����{�Sg�Q��C�5���љ��:n�sk�ww$�a�@����3ɾG).�z��q�a�Q?Ǥϐ1�U�v��vk~,��$�{
��Z톱	��ѣn��"�k�g��}���Ӟ���2zϪS��Qj���K����Ux/qj�e�X ��r��}t�X�j��Ā�ņ�a'}��gT��BJ־�D0�;R�6�W�[-�jSm�bĩ��pbg|�'q��`uj�����(B���˅�R�c`M��{��a�
�7���~�FP��%-��s�xm�Hu��7���k���K�C0�^�&C$Պ�L���򍣱&�]4��²������_�]Ƶ��cɀ��P��ʶvv���ع�� DK��/.a�ۈ�6(��<*�J�e�4��^G�|��q��zȵ�<��5����c�{�5�`{#�+���r�y�Dᙞ�8d��q2�li����m�NV��d�����X��`k�Y�^���&PJ��RIV�6�1�3LC׻���IYJ�tZ�`���@�+Y���_�.�O��dd@BK��vH%6����@�2��W9-�3l��� 4��_��0R,+)�x7��_\]�8ޔ�x�Ꝩ��K��Ir��i��uZ�m�)�Gh�w��:pN��K�f�u�;@tr��
U�ݢ��Q��� ��E/���7D~�ᯌ(z	i�^���^	`�@������I��3\����!����iD�C@�K�2��"��xrG���o��}B)%�o�zX/��r0og��0�K�n(�,�pm����g�"�켴a�$��Z ��Xз�k!�n��z!n�/����3��c��%��Bl^����	�bb�;�G6��3���T��@��u�� �Mx0@�;+A/>�3�y�#��=x����&}��N��5T\L;�#<��(����'=H�����k���.�L�ܴ�:2n��
%�R�r�����Z�xa�F?�r�{~w�)�P��L'<)_4�U+�tP�G����-n]У�rW�Y7Ll�7��ʊ'.G�{�Ld˓�����
K4��Չ$H�c��K>�\���l/-�?���u/��
�:��C�H���3�>H6��Ǯ�VE����F��C�Uˊ�D G��L�o�8H�v��b��Rgn���A�1� ����Q"�ȨÃܧ^=��۾�xP�<�/�#��dO�9n�L����#%�o�l��(����� ���=�����������m�쐀+;4Q��[���8��3����Y3��?��2���͚N�C�)�>� �`���]k����ZH�udh����Xb˓���{�}ϟ�z�wl� ���������t˔i
�*.��p�
x�HpOE���⿮��=[�ܑ��t��)%����#��w���zօ�i���&������W�g
iG�^J�xG_"�E���S[w !��I8���vq*�R'|�1]����'&Z�SP�M��Z����i��)��H8�I(�q��&��z����Lf��\�7%�s�($b��s��C`Z�D��/���ؒ>��-2�~�ő̬9uT�q��IQ׆��3�p�h1F{�>c7ǵ��T�(	N9c��ix&r��eg���6�/�2!�LZ772��]�ղy��Ց#W6�U���O��DH(坝��Mĵ��Q�'@
>���6"%�Vc�"gtq�˻r��Uo�JR��>������iwQN�i�zwÈ��~��k�d��,o�: i?�x�X�x�����7&�FNk����m7�#���s���$@k��/o:˟�H�v���ӆ%�����"b���S=��� NO�<���g�v���7+x���Ɲ��������
t�v�
&��	����:_lB2;=�o�$�^�yb�I����^)�ڮa���ߘ�G\ŢH���d�+�@�la_��\Tq�g��hMu��;�
%!`lFu3:��A�>	�r���<J����Z$��3���R�	p ��Xs�3 �[%?�����$�c|o����v���jw��lE|�2�&�	s����5��+~�3{���6��,�&�c)m��lI�M��i�o�	|�|�6��H-C� Y 6f�ٽ����"`z�=�u��u���s��ʹ���7܉T�����M�و�OL�8��+�=9��U��<��7����''b��Um�F�r���g5c��r�� ����a�?p�6��&\
/=TU'J���Gm��;����|�	%��xsB�� �W.j�=&��j��f�4�^+(���2ɠW*�R��V�"lWd����z��w��=��L�a�y"��O�*ʎ�Tw�&����� ���8�^I!�ߞV�xr�7�Y�z0u��^d97:�h1;w5Nԗ�LM�D$vq�W�>$��H�I�I5 :GFr�����r��^q/���S6�*`Nfբ��%�f��F�'
�ϔ��4VRwD��O�b��9XJ����d��⪃��-�?O��������б/�'�]�����X���k��85��gk�;a�-�n�K�IӍ3���'͔ل�Y:�2������d�U[%`�|������1Z�ߩ��Y�ڱ���Z'��+��2(Y*vn��Z�N�)i�P��sʏ.�&��֬�{��H��R/Z��%b�S�c�5��l�2�?��<�Y\7����;�-x�؅A���G ���m^��+��/p�DI�q��k�p%�������������H(Bq��6$��pv����r,�$3��ڌ�������gϰ8g�����ʖ��c��-G�X���lN��࿼"�J~8;���_�X@X�n	�
�']���*�t�L��N���c��g��A�&�d�
R��Q�[~���O`Ulj^� ��ļ�6��<vO�:��j�qA@�D�-�L�).,-$ɴ's��Hn��Z���8Ĳ�vU('��:�mՃ��D���"��."lO��&�u�l���]u}���
�+.�CȭR�A	g���)����pC<�#j�����Uh��U'�o"������f�u����,���0�_��z�¦j���A\�<�q�c�+�zp=���-�s�3��>������8�܋����r�:�'��W���)��-p�}Bg���TW%�W�˘�2�Xq��o�dpyr�pf����K���"���I���6�z=��5��ii�i�ݸKɌ��.R�"�ۧ|I��u�d�"v�����؝����Ď0�n�V�Oi ��)YsU�� h$W�.E��7�ҋ(H�C�v��ц�h�������$Y���V�W���r�� �o�����x�Fk��o�L�\6<i�GJ8@[F���aOG�}�A٪ێ�s�W��#j�u��=3;?�W��_=uk�����m�,V|���(�������H�A�7�_|Sc?�\Q�B��2���5o~�-8*��]m��e�=��=.�E��ܩn"]E��f���๊ʬ�����UbJ���)LJ�RTF����c*���p�_�D����d���f_[����Ҙux�A��z͆��浴�*��P���쯚0�%�ָ�;D�F�^������5q��㵱�$�q��aa'� ���T`q2�
:����gs�������ē(�6!���a}�p�#�n ;�/S���~�Q��/��� #US871��Dz�MsI׍'M��Z�Gگd)`�K�Vq4�AO��v9O�hB]^j�&��R�M��+*U�"F����`5(5l>�5��:�UW�;k{�҈l킡�1��Ҟ��]�n�<*VГ�`D����;�7U�8a�KJ|�Ԝ=���������)�)��^uTN�CY��v3G�|��("����y�~I1�T��X��bfF_�tnh�.AyC�n>M��,�Jjf ��-X'��_Z���ֆK�%=+�T3ʦWIB�|)aesºq�Vٻ�p�t���C�{s�Vk#B�t橒�)��?�͢�"���s~+�Y�`,QvR��0.�`�UQ��c��|�n�=y��Z#ܶƕp���f�w��+jO��_q�AO��,|�Ck7������P?�>]�߄D�w�Ҋ���M��kLo�8��GB\Fq�D!���`��)"�^?j�s+�MŸ�z��T� ��0�͋?���1M�EXd?���^��d���m�Ҽx�������s�M!ZuqQ�mX ����m������b'�^$�;�9�"^]"@�%���4?{���v^����C+%-�+4�vW�n{�op
N�rh�{�D3a������+��o�y�-ىmQ�T8�>q�����i�����r�#Q�9ڍ��|wy t�x�h�09Mo��5<f��?�2܇u~[���G���a})��#A����^�Y���v����o3Z��7HN�r{4d���Ԫ��T���z��"��n��vh���@s�W���[ �s��ҙ�TC.��ڎ�7Ce_<��w��R�T/�iI%W�R�Me_�`�Q�
_�Hg����WƉ���}\�y�}6�;�ѣZ���v�!Gr���P�B�HX�������ޢV<�f��� @?�m�@�^W�`���leq�ԛ���`� �b��`�!� 5���G�Ж*"�iC�,��м��ŔL�ǟ�i�Kg9�R��(���_�7�b:��w�[�\��Ѽ+�B�dίtKȦй�"��P4<wg<[T�͠4d��P� ~ qj�Y:!ck�C�����q}���ԙ�k{W!�LB�x���Kw�r�n���D�H�$9%P���TD�30�N5���r.��!�j�k�#xZ��-[���;���\���x�jgq��� �L{df� 5A]����>o�B�+z =��7� �c���'��m� �M�5a��ׯU�޶�'^Uz0T��Bw9��0���#U�h����nq���}(�ɗ�2��U����$*� m�&X�Y�=�r�nx�_��f�G�&�O P�-o��V&��wS(�s4P\��y�4dK~\���u͑fs�����D�6)F��joO�Fփ�R�1LK��b�1�*��Ӥ:a�<,9����]�i�ځ< ,=?x�ЍJ�����:�{����!���;��;�kr����V/2�e�$�(�~���_�����^��|���@�5}�R�5���#�������F|���B'���׃��U`K$d��NS����l��_�o���%�S9`�ݢԄ��u+c�|��}/F[�'T*�wLZM�2˔֯�)$���Q�;ʸ_�j9���_�E�7"�������A���_]#�v�@�1����W��f�`LF7Mt;y>}�Wlv���Xd4� p6Ƥ �2�x+@c�� /Q"F?@eOB��G�[x�>� 5Q_k�iz�|��<�v�ѹ��δX�u3/a���\Z5�߷Q�Ŏ��Q�����a���\�e�w�C��!�~�В���/6�#=A�_`���S�7��][�@�z���P�5�K����;�ID���8��̢��@�g�+�t����\�P�����#8ĥm4�`�c�A�ʓ8�@eA���*���J�
�o�ד,�<In�3����V��*9MBt"��1ǣ�R��r �����h5���0�;��#|A��	w����޳X�~�R1�� ����Z�>{7�%�+�:#H�zs�$�?�44��('j��P�|��LV!��G!ވ���Cq�e9q�&�@ҙ�bӁ�|m����Q)-�������]6�m5�8��1�zR"7�B �ǭP?�^T��V����7��O-BݗiE��'"Vg居lևZ��.a�y�H������ݗy%-�*䉝�wU6���;�o�KX?�;
���
Gt���;�I1{w��� �y�EWm�Ի�#iB��X�D���/U�@���k�����E>mwc���ω4��<298E���D��T^p.��� ��Dl�y���qr���N��.�NNvH�v�
:���xG�	E
��{n��Ғ�I�U55c؊�Ծ���A���g�b�`�W�4�23ɝ+�'1���jG���9R�]\~�/&ô��A�h�ƻ�*7�X�z�h�:Q�:�Xɾ�ǅ�(��	�"@6 V6��1�H�Oǡ�jTE5f���/���1~s�)FS��`��N
��YfPKXR�p%��F]�`����e�/Qj//\�R�`U�c�j@'Â���м����p"��Hv`/�[��T���$�S�'~��>��+��㥞�<X��֚@�L�ߛ$B��j�QJL�+�K�AE&�+�3���Np��y6Y��U�G1L���`����Fh*؛��{����Q�eO�Q�$��%y�Z4���ryΕ#<m�m �^���,WR�/�)�����t8��t9��q���l�~H�+�Y���j�_�K��`�62%���3�<�צ�_ƊuF�2:�.T�7�5�%2��\����?�ZL�u� �𮢜dL�3q���u�t�3�t��h-��mx�8�{6�W��v_�sQ��3"k�=�M�p�Pwt̏$]�+e��5|^
�n,�A��n8�:L����jo%��
��6�2G ��6�����@|��a�-����X<gݛa 6���8���z��Z>�,挻�����h^EY�F�2u�h���k��֦c�-�p:_9�"����l&�C�(7NU��Z��P�Me:-��[�k����$K!{]����^�<t]!�P�*6b���YH����wL���خ�(���@��=7��D�p�f��/��U��U�k�9�������H��V��
R�B	��d'K��<}����/����E��t���
�Mف�i��]c������	z����dutᒆ"YN�?9���콽NpXRD6tFxH�������5�@y�Ȯ 7#�¢�Kw!�&$� M�w���;��2Ҿ��Z���#
��f��c^Pi�[�д�d^{�#�V��/�*��6��r��`G�G
�}k'���8#���~_r~�PP�Ԕt�c*���JF�a7�ݥ1�?�@�R_��j|=�pZx�7�׋��Ն
�xK'�"��,�}{-�~��-��i���?��л̂ �=c9�|��Y���h��J��:��t&�D� ��t���X�N�H}i���D�d���׋i.��a���!91�o���ɤ��m%e%h�e�b�[�y��n�Z)&��J�ky:���.eR�a7��ǘ�w�w`͇%�ӯY
}��=/�Cn���烞Rm�Y xs�����o� �rO������Ep�Ԑ�4*���;�g��7S$F�~>f����*�-3�'�����Ӟ��E�[���X��I4�`2*�[-!5حt�����G%�ޢ*�a�iX���*�=�Ƒ� �R���h�j������V��$�4k-	� �� )՟�����zE^#?	?�_���[�l�cOxÐ��Q�B��@����Θ�H�0��U��~��w$&XZ�����G.v�J
������n��@��Qt��;<�~���÷N}��5Ї�dd��ðE�y�i�gΈ��꼂�T��Ú��^�C��d�r�La�y�Â2���\T䄺c
����PX�V7��ʟ�}��:)	�BQ�uj/4r�X��g#_3|Q)C[dH��Yoy�Z��k`iO)2�ܹ�5�O댰Lc�:U�AR���u/=�`���H�KQ@�1Im>�J�f�
 *��	kد��xB�k��]�Q���)�
��:2�'S!��z�z��=ۑ8��;|&�6�+��u�'��أ��������3��3?�S�b�Ψ	�b{*�g*�M�9��'��I��K<�َ,��)|�����&3���S�dX�L=S�D�<-��< �(|��S
7ȃJN^�����Sc&� �So҉�D�lSH�X ��Jgo��!�hޣ�?�� �巛xo匫o� �߮�-��.s�l N��ɯ�i��ӏ8aʪ�;_��G�'9ˣ݅��^�A�ki�� ���~#�n\[]ep2j��EP`�I��[0^D��J���e*~-�)�]�+���̇y�Ꞔ9� �&��M̀Wf��+�le�4ϟ���0���d��NLF��(
 ���	�GzNW�;��aT�
�5���������n�(��f��]��hD�����T?�l>�L����,��0Xo�[p':m��ŵZ���3��o���QL@IW���T�T�O"�"K�g�۩�D�%9rע��+�hQ�٦� [�Iu��	�/.�߮�� L�q>	x�\����H[u����`��m%Ƙ^���E��3m��n���ܼ6�1��f�a�A�W r��M!��*�m��seHx�[���R����Z`�}��Wx������g�p�-𵃽�X/���}��L��'N�cg�	"�ޏj'~����+����L\
ɖ�A�
���NڴM�9�wJ�M�w����s�\]E\�g��c��Bº�Fz��|&�Sȕw����s���$K,�jz�=Ӌ-�qMoN��G9k���ᾷj�����a�6O������s�yI`�(xt���X����10��$��d)�J�@Y�Y���u����
?hn�����"�鬾̏����4UK�u��n�|�mMJMVZ���d�Q�~nSx�_T��S��
�-�P9��s6D�YP��z�yS-��7�J�{Ғ��N9K+��>����C Q�l4��_Q'��(XNѾ*1�c:��>;�c����<�t��8Z?D�����eU�����"e��Zw�|��1�X����h.F�#����C ֎�Tn���|��* >>^���|u4M`=�.7�.��i\r_]�$�L�;��/�-��I��hz�S&?���Kp4�z3	m�.T���.���&0Q�f��$�3��Ł��gd(=���0t{��� ?xU�	�0R�?�:P��8'���B����K�&6+=�d|:s���{I�ǩT��z�!@�N��wj�W�t�B�w�o>�.��E�^"H-�g�	8��0�ji,���%|��l�J������L|�a�d,cC]��@(X�ҽ��m�95.O�>ǭ	P�ڰu<i����1X�Mb��6�Un[MD*q��tO�kB��!��d��W����{�����L����i�ދV\���FXz�a��G����в2�N���h��\�<���G�/]*w��Ď9Q����ȑ;�0�!��N�����.�Z�u2�Я�YYOeT$�)?,��4�<���-)Up��9��Y����L�0jB7�k'�����QW22BYѼ�ns�,a�G)���kb|�{[��s��@��m�F��~��H�ά��\V.�9ϟ���x�l\��A�KZ�<�"�X�&$�;����5��2�I�x�DV7�'��[��d��"w���8�c����C��k�����)��O
�Y���������Q X�3L����m�7�ۜl?�A\����$��2�c�އ��	�1�a �q,�v�T=:t�T4&�4G�줧)�d�LB�z��K;���^���焧���mޥ>�)��0����A<a�0~�9��ǰ������0����`��v\�^=w�����F4jߝP�7I�:$���WQ:��)��1�j\�����v�����F} �	R�?������6]N{�
��i��Ut����S|����A:��bB���V6w�˱n��}4*�`|�J��4���-�Z�7zy��|��Բ�3ɱ�S�T�
������ ^v�H6�\3�N ,\��s@M�M.���Z��E{������|�;sQ���K�MY
'�m�>�b�5H������p�(���| [7�W����B���Cw�	m���V�2��y�V�R��P�p���rUB�������n-R�ȷp%&�v��5ƻa:@�kc}��]'&OH7���Ù���8Mr{�EC8""��7�Z�m0&�{]ͬ������ݰ�������Ö��}%:�m�I!��ҥ�S�6������sV�f��GN�t���뉢Ѹ!	C���s�ԝ�̍�Q2�`L'?\�@��t,	�����7k'ީPfBU:�:t����(��'R6&Nn��&T;:ѡs ]eh�ӏ��1��#>�mu�g�B[���[}k�5R�gj5Ŋq���\K6yץ�ݮ��-p�4�5��w3�8�ہ��������ی���˒��PK���K��j��`p��>�g��a�@�2�@�_ʯ�/1%�Ĉ"�-�D�ج�R�$&�-u��a���5�oɠZd���۝�����a�yI�vS�[�{�� J��e�{ZQαg,ʜ)�.�7xo��7yb
c�B����˴�򩾰L{�BZl�Gd���q��{N���'�'Ga�F�I�>���m����89Q��r'�߲8&�K����~Npw�����~Ձ������F�Xry}P�3�e�w�!�p\���==%�{*�3�ʶ��`�5È�\�6��# ��I�����2|�V����k�x�i�t�t�͜]6Y �ӓ�����xÚ��@C>`�����%\+�:�v���(�ٓ���߁���~��>��P�:Tc6� �(̓�]�U	bY��5��ױ=�}�y��c�����t3%
�J����3��E9�=�,8���U�W���/����B��?,>��M��C��I,�§�,t��!,B�0Qʟ,�Cn�_����Is�v!��[e�C��֨.�G�J��F:��j��kmi"2���׽v���`7o�Q?n�ԫݮC�zt׍b�B�}� 7��٪��4������4�淇5v=����L�i�Ƈ��k`3<6:��7]tVө�O��hQ��k"g��֭0,e�8iVP����rJ56���!{���#8;7@��Q׆xwo+@
�,-9�!���c>��\�j��m���/Y���4x���q <�3�.�<J�5�Pj�����𺽜�f�l��v&D&�p����*������Y�]-�.����p�<�D2"�����G3GJM(��ݴk /o���hn�M_���T���T�yCY�B�S���7WRY�A>Bդ�9^w�RF�/q)�O-O�0~7��6���(Y�-��8����`�4`�w��aV��q�xu��tR����kg�:Z�e���Y,{�
b�e�χ;
M�>�۾Bp��>����p��OU7h1����͎I~� �?_2a
�]Fnz�\�n��ֆ6V#��vZ$�f���ZC�?+u���R^�6����Zi�i�� %!<�:Ő�f-�J�������B�⠔�>��ȋr	�����_~=}8�>L*�b��v�w<�`Q�����`�1)�j�7�}lA�^�L��i��?���%	|S~��-�<[ZO��T���hk0���p�}�����v�U�\)��])o=���ۖ�A^�
�R�Y�����y��8E.8u�Qs �����+lK����l}����L�V�Z��F̏`:�a�?��!����%;�r\��g�0��9��Sm��ȯ۽�gDH�s(Yj5x�&5��;�Ū�� �1Tw
������)hz���$y��K�Ϩ\W���FQk3�idՖ���-���/�ڪ��%>E?O>�ʀ�����֭Ӝ�X�6��.��Q�2#����l0������,k�2�>ξS���u5Sk��Km�&a�7�|0X~�T�"��p��z^�Kզ�UA��r�i���f g��%G�t �v���,�mCtpz��{�JCKPIl����i�}�8UΡ�f�p��Pkt���gB0�=N�@ӹ��b�����T��k
u���I9�F-�7aK<�C���b;!�j��������f�<�Q�L���Q�7�]/�A�=��_��:�l�	�3��v 6�܌��˫؈ ��6l?���XyC�U�s�:x�nޟ'�I�*�/F�l����ӹnB�z�;¤�K��e�lhS�{լ϶��ˎ�ݰe����	������~�iw��hy�k^�i1���d��Qw�c�'�G d$��ɽ�E�=��|��Օ�
�Ȧ` ޤ������Uۂ�9�l�]����Aa�g��$ˡz?=�s<�/��{�(�!�[䚖��UbA����\yi mo�,g�pI��G ��ԗ���heV�Hg|A{�W+�5��>Z�!Vmz�<�-����Ԝ`T$�e�^�x�q�"Pǵ\8LO�:���R0N¸��\�ݥnäe�N�)�Qn����+�W���٦���17u"����s��8�>�M���>U�q2$}z���%]�B"|��H�};Q�˖8X$x�R���l�G�O���A�Z�A�&�:�����(�{=�J��y�X=9�)$
X�btg���g]M�V�V��/�g&@ar�n�yU7�NF8��^J@�����b2c�_$*��^�N�q�ɓ/һ�G_��C���7�w2o�w#�����H����S�xQ1�=��{����ܪ:��xQ��$�6��G��s�nB<_������Ϟ)\o)s4�ea��C�r+�7�a>9��°������5#		j-yJ��2ݐ��;gI�B��c���V�ߤo�e>�2LOH�]��{�%@�nM7E%��1D���e��$�ic}DcQ����G{gqR�O�{��鮳̞��>���D\�����]݋D��y2^�7�`O�
�2�1g�m�u ҋ�˿mk:t���e`�|��ŖĻ��#�+��ˠU�?:![ꁝ_�:rX�M��^qV�8X�k��UƲF�s�����p�6��"e|�D,KJgԀu�8@�0�?��Z#.	���z{dh ��B�����lş�Lc7����Şn�Y2�7�X�5oY�3����i��5�5��[�wwN¢��o�)P�u�|8�#��x7���ԡ�&Mw��G�� �ՐY�v���F=ơ�ĳ��e�V��L̀:����}~o)�j�";�م�\j#����ز�,� t@�I)>�}yhv��[��coA� �В�Ѧ��/3R�L�Ո�I�ҥ�YmG�]�	�Ә��5�:�;J��W���6��U�/	-~��U����܍9�)X�`}h*�`k�������AYR�	�%=בּl.���9̱=p�+�OтN�ռv�y�h���$H%s��l� � i�R(?�KH��Kh�<aаO|���l�+Ǻ �<:��h>�"�%߃��\[W&E{����X�pI���Y��'��5^?wD����&Zf`�.2n(���;yu��"��)�&}e'���`/Ֆ�������ݨ�*Y�vٖC�T����MJ�FE,\N83bC0�>-�q��m�)��-U���2��jC�^��"�H>MRS��)�&���z�Z���Ҕ���rB�B q�E��i�ܦ��:�"_�_��?(��>氯*g�1�-�~�M�򁀬V__�';'�E'�D�k���nAu�����FC���;SW]F|Tl1�G���n�v�I��V�!*��F<��*|���!W�/�d����_�p��t�D���R�R�i���#u�[����l�����ho:�Ƭ��;8Q� ؞^��~� ��޹@�sk�I!�'��J�sW��(W����WØ��c������]���y@��zw�h�?�m�x�#.�C�5�u���*l-��a�(��fZ�����I� \"�K�{�����ly�� �����s�а�.�A�YK3���1nPox?����Ɋ��0G���ɷ��شᾃ���4����O����g�/��2��V��aӸzp��y´7!�����8���@^�{�9��Y[�5m=-�8���s����K�d>&�����J;��BjUQ,=��.[�����e�SϏ�/r��N�����J�w~��WZ����1y�j��U>,i��[�s��^�k�V��uA��3������3]Wb��s&H|๺��\r<�uab�a�>D[o��8��9�d����Z�F �N�4� ���/�ɿ�0�ܱ�TvRy�}I)\�)���#�EL�<F:�},�kE(�^�'M���a~���2JV�Q� �ei��4X�> ��*Ϧ�}�����?L��n��j�$KB� T� �^s��ޑ��;������ḭ�昢������~F|.�B�����\e��EC\�qY�._�֖��������:��������2IkH�����n�Ȁҋ]�o���R[��^�9�Ƈ�rv��9{�hx���|��It�r�B��m����y]2�>�������u�a�p�>�RMnsDX���zqƒ�!7k��)˘�Q0��>{8��Z/�1I;,��Fi,G�o��q,����j�L�iS)�׵��j����D���bы��q6!�XiJ*I���ٲ�y�R���-�yAp���Sr��b�e���O �C3���Qo5.�7Ƿ��t����@����LO75��o�y�100���wT!��K=��>���]YX.�z6�5��{|�V�E����6�ބ,��GX���aVzYqE�*��j����ԠaCѬ�t��iӏi/�X.��S����m�ɖ�]҇�����+����|0��Fy^Ԩ<`j���`���5�D�{���	v�^d���l�����	�B�{�x��_�J�?q��� 6S��3�!����E5Vz�OQ�S��/xT���?���e'�)����,�~g7Zj�@�g���3.�`�l�V/R��j���]��O����947E	.�H��f�e�{C�c�M��eQ��{��h��q����Fװg���=�i�o�a�u��K��*4�ΰ�m����}��H��H��ɕ�*��O
<�X�'-���:e�d>�f�k=�dzY��;�4�9��@�~I�+ 8P�`�����I_:�o�&��z�_����Uc�@�M��,�M�c�^U��H'�E�k�>8 g��Dr�oz��:�B� ����D%@����r�.Ք��6�\���A:oe���% à� ����o�8���_67�+3 2ET��<��]��f�Ʈdj��Ա��?��'�*D9�{�Q9�fLq��w���	�OYu��=��9��e�*�N�Q��512���6�N|Ҳ�D	�\�i���OC:s+R���_"� �0q�kLȜfO���c�m�H�Nlk��]��܊9�$�^`+�DW;Gy8����\	>���=	}�$����G��Yo�A�_:�,�MKg"���$���'��p�=�l�$`/���L�.ӗ�X����JN/V+O5�rQN�C�������,�N� UѭF�qQ�Z�?(�_Aig@¶��z[�{��h�ǆ�:�x-w�w�Q��:��>$��4��AZ%+�X��ލ�a��B�#�����F�Lt�C���[o8��I1� Y	X4PL������x�xB=�:��;O>-��ѹk������\9	jEs�Eҟ[�q�t9[�����
��:��xˎ�32���F�l�D���&0�W`�#��G��b�_��f�����Ǵ�k��#���aˠ��᧮>��Y-Z&U8�������ʺe�Fb4v������� ����M(G�B!�.s]�����q��������_N� ����d�j�B�����۳�0�C#��()k�ܒ������[�-�x�$��U���ƴ�@0<�qX���|S��;k!k�M��r��j���dF伒�� W��XA�)h�\AP�����2��M+.�,��+��/{�"��3m�"M{�����F���:U�49�g��?�wp��G�R����3� /��]�a�p5[uV��y�$����U2�]���C�����^me%㪀���<O�7�E#Z�
���E�'�~�<�Nhs��t�<,F��yw`�<�! ey9FD�H0W��quHk�nj��ܝ:�e���CA���j\�(8/���زDnc]���z3�DJcd�w��]��P��j�a�C����������M�Le�بO}\��_�U[�6p��kh�6��5b����B�lֲP�3���ew ?�Nt�������d���%�{۪;<M�P2+�Ӊ���U��<�<��Sv��,E�Z2ST�S\{z�0XB�M�z\�J_]y�- ��d��2����!֢���G�}@���w��__z<@(}�$Y�q��&��TlP/+�H�}�T�L�u���V�����+3u�w�J�O����)�P��;�
qp�~Y��q�Y��A��T�5��'V��E>8�Hc��#�'��svf���=�qޞJ8Xv��L���^�7�h�.�.��p? ��M�O�Ilso�|��2�J����AR�,��W��A����ռ���V3���d�BK���5<���L�)+��^���{L����Nx�kjUD���~��RP�o���^C�#��M:Bdk��^��vU��OV{�MI��d]9H<� +�÷HΡu=�����$�s��X*F�&�1]L6�i{� ��
&ֈ����h���{.��jxMA�`�;A��dN�O�V�j�`��o��i�:4���NzyUj�ܼ�%��R������]��i�B����>j���Y�ޕfSi�9H��+�{v{�������8*\�iMR>��I�:������]xlH��[���h!�^�������.!�ʲL�+[]�~��V /��<���mI`���Jف%d���4�~��)�oc�Ѥ�J;�È��C���M�G
_R���:���_��Jj��
�q�c9g�5=w�Ijfs�j@�70�lVI#uƘF`�藓�lJjϺ2�9�g2X�%�Sȕ�-��:���ж��\c7+�R�7n{4�m�ť�UL�vc�.0��w�=_���t�o���g��������)�OT��M�y����|��Ee[�������d���jƉ��_E���W�c���:�%�M!��.~_�L���y}�K�ʑ�f��2��z.[��0L��T��K�}dJJp[�LB�I��P�uC�~�����>܊���j��bZq��D2k�7-���x��m(��?�r��}���6���5�뾎e5濊Jn�g½����i�tQ*���z&5՘��r^9�2: �;�n��K��-�u�0>ƺb=��i� a�:Ӓ�KZ��+�Ioܠ����(��7���� �����t�IjQ�q�F�N�n��|;7wH<�Zx�o1Jvگ���Q���Ȋ������2$dj'�M�,!Ȅ8�hR���M����n�Z���9��e�-)Jt|t9o�F� "���`x�T�ܭZb��-������q�B�\����(��U8��[�q�5D��b0b���	[\�C�{}���bq�6��TD-�WI/�2;��&���
���������,Z!�4{��ӑ��vt��|f�bQw��^?U�n�U�b\*=ɍ�e��-SP��+����.#N�*��a�"-m�_��`�*�o=w?S�h��3�|�8R
��38^xo|����_2.-A�
��c�HsѺ����;�1�MQ�yT,�#�A�d�Qv�ki�`2Wp��b��:N?9'[&n���$o�g�7 S=>�S��s��������z`�o��X��Hf
�X��, ڿ������q���m����ć3~MOA�?��uYv�"����|��[����g9"�G}�B�L��_�5�hXjD��&�^)��1��5I.\�{H-�D�6_�;�P���ͼ
��U%����Z�|�3n���Ⱥ����PX������N<�2&�H�j����?+�ddܭ��R�|.�
ހKB�ܳ�K�!�Rk�����Y��P�4r#�흩>FO��Hm� ��]������y��) ^��}I|V��r�Y��Ʋ4m�0�O�.:��/�.�{��O���{�QOYu"��q�>:���ܝ-""��˿��5R�w�[* ��ꂭ�unΛ^S����s�0#���߭yLZ�
_mV�BҔ��ˊ�D.F�<Ս6�l�g������K�iH�l�fKb��5E�xz]�����W�d��^����4{�`_�a���H�d���w��-*(����"�YC��)B���-!��Av�$��"���68}���d8�0g�Tf*��iL��O-�l����*� �=\dZLM�{E L%~��[.�)�K�M�o�\�Jᤔ��0�.��6rq�^0�d�����w�\B#���^|�/JZJI��5�x�$�i�{,&b�l�4A�g�Rqg�n1.;]�����A%\���"4�F�NU��'_��0г֌|��85n|� �O�O1�n�2[X�eq�f�{�#���$�%P�BoK/�<V�L0.҅U�V��X^�<{��BS���O]�
�}�K*n6v�q���z������{o�Q��&>��%�>;����%p�� �=$�ʩ�SC�_xpy@��;,��=��Q��c����h����~�GX�J�wMi;�EwA������X��\�2��� ����kx��\�	�qM>�s%7����ʖzE���w��p���%�P��V��Z2�)yX5l)`k܋���Ag-i�Q�!��X���|�	�߿H�?�"���%�R���*�����NJ�a�[�^p��=Q� ���{:[�`Y��-9��{��K����	�9)@�h�l�@��.8��h�r���Z[��ɇ`�x.߰�CN�W]�8��+�T(�������=��b)�z��[�d�L�!�_)A&����kNS���I�*�"9Ǵ���3��k���I]�%6�u=��t�������[��8�b-��xǾ�)��dC5����6�2j�IQ����`��)W`ʀ��R���K-,�(��� n1��j�ǩ�D�=I�ܗe�/�����/�5��G3vE��_���Fb����}n+^�LW���L���F2ЁE\o��;�t���~ӫ2��S�R��(?��:�.�JlV�jX� x8����:;��L��y�1�����[��N��u8���'R���#����?�-A3J��T*5��y��(�K��Xu�B�с-��%O�6�%[<B�|�`�)f��=�,n�04�)���`�U���A
*>��& ��5I[18L�cG^/� j��%ᅔ&QL~�C�`SY*�ݑ��N��0-�$�2���?�0d�1�)+�Y4��e�r�������-�����4�s�����H:�|��Z��U�-І��l�m�����\�"�Y��DU���T�g�p�Pa��OuC�M�0.D��\��u���a��P����_K瞿7�����G����vq�fr��(0(j�3r�}@�`�;ݛ.�-��r S�Q27��-d�Re絏�aB���bZ�����{IT4��L?M	8lf��������fA�B߲71�W�,BE��ʁFo)���U���Dl��Z�xH�*�Uwj��?q,�Ж���-Ҹ<�p��DD;����[4� ��O��$�h}J���c��}�w;��0>��|��s�7���#���Ȍi�_G�OoeA�"]3�{"��"�O?��o�m�t�*��0�H"��2T��ʑ�΁��In�׶��bjC]�x�b5��o�������hYé�*o'�<�/����/J���K��\s�,������
F\A8� �&{�Jaè�-�:mk�8�3}k�0o���͑�x�V��s�O��3j�.��h���~�2���}櫒�֘�B��#�`�bC�6KU�X��A�Z�~Z��)��-:F����c�#7;����ӟ�E������( �ӯ�xw4̊��=o�Mfw��Z���F��xM��Rp���W�Z	� ,��(yV	�0��W�$��}�ڊC�c`���V�}p>O�Fi��qn�`�HW� ʵ\�S�����OD�NU0N`}�����3F�g[�
�ò��:����`��h��a}��{���
mqy����V�e,��mġoBM� �pAP�%���^l�F ��4%RZ�u�ӝL�E��'?� @�5C�y����(/���$����3�X��+4&��ې3�?�Q�Z��}͞��oδ�)���eᢳ���l1��F1I�~�(KE��kļ2Q�ȠB��;��r�Χ���(�fe�l��Z��=?�/j(��%�K���	+�>\�V�b��δ���}��*��yA����c�������x.TX��ooܼt��_�������n֋S��B����X��(�տ�|_C��Wf���o�~ ��g��V�Ӑ,����m�F���ɻ�ɵ��5��xaD+�O0q�$w�8'���
�f-FpdM�~��\w�m����h']�xh?�I�}z����J��3U�BN\1 �}%�^W��,�*c=�9Ƴد�M#��+��0\l���4�0���҉�*��iV!��>A+�\�:s�|� X�;U�N/�<��#��k��$ZXx�^�� 7Gw{����!!u>u�;x������#o���d��r����MX�x���N�8:dē7-�̎
T�^�W˛�w�u~b��������d�ݥ�r�~�*}�J\����<۝�~0vOl��	z4�)H<0�3����a�.�>��c��D��Ӿb�b��t�H���$v+'�oY�!�x(�S�A73���Y�O	����̸� %��5�P�� #�y�N���8zH�����N�	d7�������9��䛑�yb�[��"\��ښy�<�QnThXF���l�vx�3(�)��9~�B�`ҍE6�C`����T��ÝK/�c�,b���^�6�{gq5��"��$��>��D���ҁ��>ߨ�\/xa�~୑>�8��/�a���P���-��bS�/�jy*bf3�!м�,
xn>�3���s�{c�#-ⰐB3�R\`�ܜw�쮅Pf07S�ןY��^@`�qd�}^��xhC ��V���]Nkc��������
(N�}2�5�s�@��%ui��㓕�E�-}.�뽰4���%	<ΌҭadǦ���c#��ԘoXf�O!����u.r�����6_7E�y�|t���o�&@�i^s� �h2�xL�T���m�����g@�X*˻��Z�᧢���[�m�L.yˆ�&�\��N�{)��_?W��DϺ��=�J<��E�jӈk!��6���%щ"�p2kY�/]r-���_M�;��Y[��j�l���d���%�����Q aL(��S�Ri�T��o�"TV e>�R�@�ݶg|U�����Y6-�F�/Dc ~A�X����If���Ԓ0��(��e}v{�ۡ3c��
�#�?����vެߗ��f6cy�K�΄�A��~	�����N�
5��8Mw���K��g�T"��a��c+�z�|"�*�|3���tZo��1W�ɴ���'1��ӘQ�a�zЋ�&�r^`��L	d�F��E��t$RP��t�x�:��/�/'��T�g�*���<`�}`+�\�A�O��\�C�^�I*�E^�e���F�
U}�ۂ4v��J��_*H,��ɯU�������-"��&c���	{S��0<�'��]�=Ã
7��O���椮k佊ps�#�g��ͥ�����Ŝp����Պ���.�����#�~~�*�MeC@?��|��#O�m�-��h��E1.� t���[����`ǃ#���ٸ�T��6��԰ؗ�w/�Sb�dmE��d$fZ��#�
�>�A�q���Ē;k2�aŘ�� 
���N�#C���R)I�֟§�7����"
���^r&���P͊�<��$}��GW���s��dN�5Z}6TŌjT��Q�\�v��3���t�PSEz,r���w�]FF�+�ɗ��}��㭌{�j��P땋�\�E���o��R����*#�H��E/����w	�k6��x~�<:,"�/��%tQjPDJ��=���g���7�H���k�;�I��E�P�0+6�(!�Kv�ְ|�wz�d�L����	�~a}h۟m��!��@��p�>%$��-=E���z6*yn��̘��X�P� �OߒNeد
��?�B��{E�U�J���B[,�&@RqT��֙N��^�Zo'uS��4(*�e|x�3|���P�
�Z�Ȳc|k|B�ƞ�V)�<����ĵ���_���������Nb1�� 3_�^K�AP�l�K!>NI�h�ΫcsE� E��5�ˏ��j2���c�KP�{�^�Oôi��AK7��Bb�%8�e�yS�E��҅t�lU6!�@^��KBU��RǢ�ak�Q$9̓>��P�h�kLt�/�F��ɠ31��e�rA�m�T̃hN}��_&� Ö�}�h�N1��wg,_J�E%��8�zn �M�BM��)=��t��N�2�������@�&����9�y ����׋��0lP.�i�\�ck�z�_�Pc7��hmޔ,�3��[9��z�����YܒZTkM���X�J�����ov#2��1�p��C�L�0�����j�&�Ä�$8���*�׭$�#B7zi,j1d��K�bC��A\�xP
�Ɲ�(k�K�b{��5t�l�< �k���D��?�� �m1��F�E�cT��y�{'����Ԙ��&�.��Ϗ^ �J6��d�`<�cu��qF���ט�F��M�c��+�N��g�{4����2�uk"ͱX!��h>e�_jb�fr���]E��J�.v��"���_��+T�<�xu��v�p�/��L��D�#�L�F�kW'��mN����S����M����W"�B���ٱH��ϐ�7��
�q2뜐lLe_�z�7P^V3S<T��'o��ԗ����E��9�i&���
4dr!����w��Ѹ50?��"S`�g�7��:.�P1��%�wG�g�0�/�6�ʙh.��qzz�mY���b����=�l�4؝5�as`��`p$�l��A��H[�a��E>u��X7��vq5acT���;X�D�Rє\4n!�E�pu�.g׉��6٣d��k�k��G�:I�?Y��� �=��|�Oۘ���j���J=9ZYf�����6��ߩͼ�XĐ�j�B;������>�d���ѱ���M}���Bj����-�;k����"���ob�� P>l^����<j3\Hޠ���Zة;�2�oV�9�^�}��<	)$u�{�+JJe�3{4M'w�UֳA�?���{m�Z"����*�7�^�9�jӯ����I�]{��]�S�**�3��QT�⅑��*�zZ+ԾU������&��<:~}7{� �Ɩ'���#���w{����"#�s�0R��f�w��HYb�$�����l�T	�/�a�C��k
����]i7�dr9���^[�t����(��M����	BP���� ؍W���_O�+��gT&��g�]@���mB�����g�1�����k�����V+�5��X��+l
s%~����mžy-�&䍟6X2�$�~@;X�a�ɫ�	�r?�ٙ�C�۴�Kܠv����>�:�%��{|��_h���= C�2�,���~S���#�����)�o^��?֤_�{ׂ1�}RݫY�3�grl�V�-{b�MuqZ}Y��Ŵb&�<�e_h#Pz@q,��֎����yd~�Ek���E
��|)����H�V���Ye����Kx�/K�l�S�p�,|�|7�d!'_��{�Y�Ε�n���9-�k4 H�!m�x�*���	���L]>Uqj.��Q¦
� In%Š��('��S��#w�"����/Tp-�TE��sX�[��+�1"�K����Sl@�|�ũ!`��R�'���_S��t�����	lY�I�oh@f��AY�5��P��vI��M<	F��]<�\N�у6 e�|c�-�J�����Ʌ@+B����ޘe7J����'=�6�Y����F9M��<fs��:����\�� �R���H�ƫ�K/�8+l�g��@o#��c��:NPp+�߮��ƙlGXQJ�;p̳�Y_*�D���P��d�f}y�#|$���R��69(h@��U$�k.>	� ލsE�'��촲��)�>W��D�	x3o�7!�B�88�F1�zd�C��\#����J?H��vڔ(�,�%rKǎ�@ �h5�p������"��%�4Gv+g��G�Ҋg�E�Z8"Q��\7�<�d�,�Hj��&�@��!E��7C]j�2�ϵە���qι���2K����uy�|Q�}�`�_�B�����N�����[����Yo��F M�kCK<�k���PX��xg�b.4���p_L�0��c���ɽ��U��pw���ؚ�nQ�@�<7�u8�Q�S������/���� z(5���$��0q������eZ-���y��[x�Nj:��|�딾��<=B:���.��0���BL����U�/�;�0���x��[���s�4������[ކm�l~�'jLE\ ��C�t��>6��XB����u�a�
�	�H�K2E�m��H�����dp�6r<��!�w�](�m�-l����6�^��t���9q�`	g����^�I,���m 	M	�!"Ϗbޘ��v�4+H���!����Btf� M�;�`|(B��D���!���(��lF�Hc��T�dR}uiDÈ�jR�n��ؖ�.Y5�����pv�!��y��t���B����'�D
��Iױ�#$Q�	. �I՞883mu�*|b%�I.�2/B>�{@0���~�M��<���n��l��c@m;k`��P���,�34���?��bY6���p)�D�+����Ex�{U�\/���O��4�}*M����j�Zʘ�o{�B�e���b���wI�B��+)���آ412�9N�.��+hp�į�	��G~;���8��<��6��
:􆿜��^�u@��b���W��u�	k�x�2H>�����%<�@R�Y�6����3O�"�~��AlH����//nɞ)�#hK�}�G4����)�0Few�9�����C���_���T%{�y�Fo��zn�=�j\ G�v۬BVآ��-7�(y��`�Gj��JǞ]�[2����H�1�  ��Ulg2wG3r�� �`!2���uLƊ�QI�����d�,'g�gϗ'��e�"�-�[5d"�6?�8X���-��9�v�ĳ}*0j�SC�O=�����c~��4�l��՟C�Q`�9��F�i.�w�σ�0�g�k⬣X&~׳daA�y�d`S��$�]�z}�t�!��Q(G����W��A[Kt�}]�3ߐ��:��m��68�Ƚ���.����VD��}k��=�a5�`,�5��"�)��O)�J��)�\������.$K�D*ޜx[����J��Y�ѿK(�<�}�
kwW�9����Δ����e��'�̬�+����)�w���]{���O_u��O����a��魈��u������#%c�4R��D��l���F��:m�=�~��k��G0���P�jʿ�!�7��uI=�l}b��	��n/�ʛ��d����#�~H�zz��b�����"�𑲫C��3���m�pa����_�+�6s��%�#����e7�Q�\�[���U�k"�R1c��<P+��~QX
�`m�Z)�FV�V��F�"f8���<ȥV���� ��2|B�!�$������
7?v��K�D`VfM��4����� w_	ř2~��o��&��Ps�%��d礪��h��]����./)I�Z&�~�dvOZ�� ��
8����P���6ɮ񣀄�.��lk�2�b�qUf���es�o���{,� ���u��b���o�BXq �9sRS|/ˀ[4�K|K��6�:"�Y�"9C5H��z�l�����<�G���z,5� ?*ä��A�g�nV����HPa᪻�p����MUV�c��IC__��̸;����"���U/���h ��&.d`����~y�6�>�6Vr�u?�V8
:���#.��u�񅷕��b�8�Y/�h�s/��X�S����k��c���K��U�$%p)��,�]�Eu�[oCWb�!]>��d�|�-�ibggL������	hq�IYh��XE��#VWf��I��(�}Ŗ`���[�nl`��hY])�<b�3�����.�w�>(	���J�e�m8�|���=�Fqx�� ,M�W���o��q�I1���h�����'���P�A����{߶]>�#����{�n1vRTRp��W>F�T��Mv��5�^�PS�Ϸ EG���M2����#�\潈�mcЀ��es��3l$��H�;���\����C*�/�`���2O��)�S���@ �����E5��R醔�S���`HO�p��:�
N������a��z��}�y�xR��e�����s6C�0�#I��E�`�5��h�,��GD�*@���ja���E�D�ΛXp��B�Ly�=v��Ѱ�j�U�|�� �<:�?:�k!務��B��*��A�8׏
�K�P���u	;�x\}/����� ��_�(���R_��{~��rR[���-�۲<�M�����2h�,��5�M��Y>7��U��l�|��){]��t&�ߣV��Ͽ���d"�p�[����#���0`'%�z{~��h5P�Χn�Ί��ܔ�f��k-���YA�7�w$w�k�3��>p��J\�������}�Ҽ�3"��?κyò�*�נc���<����L��	y��i����m�
�[-w��]|R����h���p�|���7S�C]�}Ou�4��Z��P1O��MP�oR[�yJ@�Ջ`�z�
x��v(b�����;Wݶ����RCJ
�B��z�\�p�W�iÔ�aMI�P�2h�ǘ׸,.	�E���p�������/��������I�i�Cm�#���6<ejO�b�&����-}�k�X9�$�c|M��<��&�����d�@:�@�> ��6Z�렫f�����k�씴zj���"���z��<%���T�$�W�\TwM����Y�X�H%�-�C��ܢ����� ��+��Ǚ�_}\/sk�5��}O�M��,�!�t��<6:��%9c�i�)�3!�s���8?�^ � �K��Ž<}�s�u��fpp=čWP�wi�V�=��&h�^��'j��7l����If��c�?<�~�@���"���8�dD�_c�нH�"��8���BNI�I�N�;�hҔQ�#	$'�_K��>�����=.���,� ��޽�#��3Y���������k��'H&��T)�,��-z�V�H}�&{��V�b�����d&�������$�a5I'�޲��L��֓��su_���=��rΔd�蹘3Ƨ�m� �`�C��:lf?�ck �܏|K��e�I����/J���8��)'S���WN��%0y��'�q<!��&'���rj�K� [�p���[�Ѥӝd����;�o؀�ul�ÿ&��>�z`!��)���'3��%���ɯ͉1,�3���lr6��Arp��!7���o�6Q��m���&��S�ķ;�q�|ma[q�WC#ջ&�������U6�l��x��oר)����4:r�a���d[|�?�-l O����	(q��a����~d_5v�0�U�0�)|�f�M�+��8L��_�V�+�� �<�{�[�l���8�w�D��$1P`7��!��:����ݕ�!�- �<*�V�Y M�w��f{�������Vj�Y�e��F�ذy����∈-Қݤg���Q{{$E�뷇׊���2H*������Q�p�-���+��$�{��:f���ٰP������m{`;ǮW�PX�x�*N�N���-	��lg�r�X�k�� ���q���������~�#�L&��n��;{�$H+��M� ���C �b�uD��\RQ*��!A�NB�R;Wn�ز�~�����VZ�I�D,�i�l���>�f��	l�n��R �c�x,��gzLh��JR�����W������d}w�T�%�g�T�~�p �ЀV���Y`�k�M�c��ᖄY_u>�p0�I_I��}T*6�J�������S�?��Λ�7_f]R�hzy�+2?"��1N6�٠�{{�9sd�p�K޳͒N;Ğ�t0�
�����D=,���AE�>W�Ǔ���Oh�P�*aVHA��<.ud9-n)�]?�y%�$Nⴰ8��;�T��Ry�n���ΝF%�hj����_�(������������{�¾��=$�m�|?7����/����'�~c�L�����T�3;�����W�u��N~혴h�*�+u���@�0�&�u��iv�t�;��6����x)���v{��F��OЬ�MP�ܭx�ǘUm��{��D�*���8\��K;{�ju-F��Lݒ�GL��٤���/P�V�5�8��zj�"Rk�=�U_�5&�\�;�%�5)M׈S�Y�Z$}���EUےbs�}M�5�\)��� 7���w&z���'M�1�0}o:������9���%r��8�_إ��_i�u���2�d+�4c�
I���;��N�hBPr�K���!��	3*v"02�<�X
��*�͎DNMڞ����ً�2~���!-V�1r�|j��?�w�)�8��il�l���.Ħ�N���TI�����n�����6� ����ٵ'����V~d!��̹d�H���0�R��4����a��J�񨂭ڊ ��ɶ���*�`Ǟ���&��C=��9-�n���E�����&-Q�dF��ã����1R
��ifBTMn1o 
�!M�83b�d"�0��M̭�	�MF e(
�kA�L�V(�bJ[)�o��}�3
�4��b�1��d��ۋ<���ز-��kF��{rERT|�����^f5������=L0���� C�B�&8� �w�.�Ʉ�]Mv�s�c�k�R����h�ۭ<��Q��z����d�*9�	��P�a�
[�I8T��J;$	�6�I���,<8�)�-0�/\�ć�\�hEJ�b��I�pX)b�1�� +�E]p�s���[0��4"�Ip�"�I+�iDxٛ̅��{K�d)���\��D�I��ypXT�����[�/=tV��=q�G�9=�?59�o6�?���]d=vw��o��_���.r{=!�/<s�R}�������X�Ϯ7�y�`|4#�̜��Y�e��i�]��
4�A�:���8�CC2�H���3��/��Я"3:���~�ّ�)���7�c��~��%�^J�����c|q�aR�|�0�����q�)e ���2�a�P���0��'��r�?}`��hƜ�h&8+y�
����i��q>B��W��Y6��]��P��:���E�Ρק�S�rTu7`�B��H��шs�����r�'�8�p���iPو�b`�d@�qT�"��
��m��MZ��R���Y|b�9N:�9ۖ�<Æ;�K7+�J�]�1b�6J�r�iQ��@����8�蚧����&�(n�Q-��G���z��#yݩ�������eb�~r�S�9!� ��̅*'�1��e��gug��0(j�g�Ub�j.T5f7>��#S�1�&}��TrJ<:���6p�LEt�r�)�'ږ���?e�*��+9;���a�q�ܔ����Z�{m0BD�}X�#&�|H����L��ӧ���9F��*�#�r��)s�{��K��t��xW �D�{+��Z��=�����v�G<d)`ތ<�̮�W �coel$r��)d���Vq#��d#�������Hm/.��)",���z�	�:YOeV;u�qɚ�aG��o����� j_c���;ʕ��b?ҥ��S"�E/bk�S���O{�l�̼K��;(^�����g�t@x�~�ĎJG*����/4gk��$�8B��'g�vƝPA��8��mv��r��ٷ�H��[ �U��)��i�Pȩ�"�r���H9�� �,�J�WO�n�#|��pDe�Z�wb�!h=U��:l�/��ʕ4���'�����Y��R��A�Zթ�B
�ڍb�o���Os�%���1/]�t��n�J=�û���|�Lj0+���P�3%k��d���s]ߌY���yQ������cPz�]�w:�:��7��"<=:��o�����	�#�9�i�I�Cɸl۠�=����[2<�PԖ�IӨ�ܛT��p�g_
S�H���0A�KN���.�T}Ji�{#�UV/rM�8�����m����Cv����7��Su�S�*{���,)κ��M���H����Q���y�?K��� Ŭ�l��rv�$f�_�G����s^+<���G`��D����aQeY�bŶ%�M8�$q�8k��ߙד����eJۭ���_P���=ݧ�������s9�� ��V��h=/��Y�pf6fFd*�v���"Rt���J{o��6O��p=({�Q)��x�+!�s�I��:fr�ª��8�U��xb>'�V@Vo�)x]����j/v�?�1����+�.O��̠�[k*�N�-���6|΂i�}K`l�M�|i5k���A��.؀k<S3���U(��QӜɭ�)��nt��6̕㘨��`.��b/w�<�������&�+.�z����z6X!���,r�s��-5b�O;�cJ<��fQǚAq8��g������W��$����z�o�#|�}L}{ФtT$D.w�-����䙮{�,ațl���`�� �=
�t_���΂6�	E<��
��w��p�id���F·r��N;5���"3�o�b���ꯤ�{է���*�ec�[���Q��+�@����o,�tD���L���d��8!<�9L����(�]}W	�%��?�t2<�W��X,��8�
�<aR������+�Ϫ�Jj��TA�)��_����/Dt&+6�>[1����
�5<Km��w���i���B����R9ٖ�����<��7�ъg.0m"�y��0g�ͱ����%�x�n�&�ܒ�[e�>��P���ѯ
�/�*s��ey�$��K+����k�}۠��`�kH���W��3wT��|�Ƶ��yl��u��j#�dggé�;Smj���=�ʄ�Y�
��+��Ѝ�Џ�: ��6�E�Tq�&��AV��Kg���Y�e�e<������@��^\��t���"
3F�vzdٻ!d�
x�U��p6֩*J�c��gL�;6�6�~ �r�PG�H�$�϶��@n����������(.Hd�p�-j]�6�X�v�D�pb���]:u�n�"R�>�;i�O-r�z�6�Ԑ�%Xf�zYZ����"b�\y�1{eZ��R�C�{[�O��qiυ���2:n�q;��АO�}�o�����Ɂe�����'�i��}�f#�'����J�R$3R�uU�L��A��3�>��	Fp���堨���q���j�i��4��t���x<$�c�#Vs�X��cDȌ��dpO/]�g������f���?e�=F�<xDŭ6#LՂ\�����!���䏋��&دO�����(w:X4�NMM���-�����[R_�oB�m��D��X9���g���4.�T�JV��h��ʖ@K��j]�=�C�����%�B��b�Z-�,\H���#��D�����Ɏ�*�#\  �e6��֨�7M�C����p��rZ௨� �.��V�KO�9���K���O�)�ʶ}�!A]�)��[R�8C�XL��]���[����*�� �T�ݬp�E���mH�t�e���+�g��q������]5F��<{Y�f��`�gb��=�����M�+	��^|v_:��]��*=^]������̓Ly��͚
��T��7K���S�������
V�S+�{O���PW�2G�Li�m��ܖ*��%|�m�~�^�QD�[;��o9��̻\��$��H!����ޮ��yj�D%�D�S�S!H*) �6E]�0d�\��<"�D-xX�0A��f�e�S�C�h?v�3ݰ���4S;k�W���R�kL9�T��ܩ���y��.uMh�� [���:��^�zO�8���̄��&��ch�u�l|$g��V1�pO�c��k���_9�%D��ߓ��w��j|�!�(�!ɥK�]@ d9���a�O���Q2�0�b��g ��o�?~��N�[=����6�B�i��[:�څt8&�햊!e(.l��i����/]����$1�I���Sx��25^u���<9��5[�1�'�7�C�s��.L��܉C%���h��g�w�z�-�{�Ȃ�
��1�	�7e�Ku���W�&��}�	�%�9T\R��F�D�E�e//^�$��-���r��:����nr���czW\M�����)WفIx�1&���2C<�U\�ϛ���I��3=�C�}ϕ"+�U��
�0c��D��;?E��}^�[�zS툆xrO�i�W*�[���j.�.��eL$>���[�}�ػ@��%	ta�I�5҈�+g9�~��(k"�"huQ/�K=�9�4 )�l�ɱ�{����.�%�z�<�(�>�_.Xm�<�a%�*-�6�Hx~��(�ӥ�z=�*�[ڲQk/ha`�U��V�� ������X�2(�~�0Wz;_tW�`���#���ZI�Ĺ� ��Z+y����
�C\��OOk3ɖa^׷���܀=����;��n�~��> �@�j�(a�}a1�*fP0�^�a�!���6fRv`|*��MG]
��_��HΔ"�;��n���NΪ�m�xdx7_���# N΄(�]���8
cIʫ�������H��	#��$ #�|�`��֮ȡ��0�݅��������$��v��u������5Л��k{p?�WPYΡ@��G	�7>�j�8VuIS$����|yI��Kǒ��R,�}z��XG��J��XR$�𜵇�~�e����ЛAs$��ش��#䷸�����4O�>(���X��
�6R��<��/�H噔�x�vD^��F�J�R��~!%W��VIzvJ����6?�<$�wB^%��%׾}�_b!djg�W*Ȅ���^��M�[������o@�e�Y>�f��J�4��Q��+,�?�.D/��.�7g+�C��r3���Y�m���u���F�t���O�˺h!=�����
��x$�<��Ǿ]p\�������8���j��6d-�yIC�e�nA4N��&P)�ȖQvf��ꞧR�|����H�6c��i�DG��yZ�G]`ؤb �N��,�}q1����X-���/l˷��U�[Q_W	��F�~���r�v��p�L�+�������Y�rx����58��^T�2����o��)y����id���w�U�ݻ,��������)�zE8ۗl�'h`�'�V�-PE���
K}5y�n �N+lrs:��8�+0�}a�ף��@�R\�÷�y�Fy����י��e��nWA��q$2�tn���P����al��P4L>�0K����5���5���p�ɿ��nO�K��bħB����[�h�)A�m���a�Q|=�����{�@NIQg����imA׎R�/؂��;����S�`��ka[�P����樠���ʭ���	H���e(W=�r���<�?�����2REh	|������ɮ�r���K�vɶ�E)��3���jU ��♀8CGc?kg�s��V�܌�a��AK�ǚ~�~�����b�!*K��o����k�#A]��sc�ಪ O5��J`60:^A����(����]��/�,�#�4����ﱻ*³�塉z�}��ﳪ�&�ɸOOהM�i�w�u�Y�ӏ���:�HD�.VZנ��6��CO����	~�T��3:A��#�-��'�a��4뒁��zX&%p�-Ǫ�Y�' �T���t���/[���P}ꈭ�1�O_BvC�{Ó�]Վ�!�ŸG��GK[,������Didc|����1�z��&	p�BŮ����҉ƫn���J�%��#��b�v���Q<�5ֹ�z�T������9ٽ��Ӹ�W��³3�^?��"[t�YO��������)p80����{%������RP�֦j�n~����6^h��c�N��֤ZT#A�
���!���"�>��k�n>6�1���CW��p9�X�,�3l�W�Rى!�����\%�;��a���������7_e}��,y��FÆ��V����y� �<z�0U�lj�e;O���=��Z������N�S�o|�H�$DzaH������y�.�IP(�pAe�{�������!�,QA�Q̗����'�ޠ��KY�UX 6�X��K�3�g���U�6F�=���6J�ϛ*�(�3о�:M;�9���>�Gi�!r�E����Hб�Ka�7�E4��|���B�E;䫼�O�=�'��	��&�u�L���J
I�[I�C*i��%G���t)�H�ۥ���sc)�1zrQ��n���Q�k��4��X�ɀ�YQ�̀�õ-��#bN����C��P�w�� �Y�)�\�>/7@h����wjY�o�W�OD�Łd�l�o�0%����u��Q�m�^G���'3ڒ����;�G�5x��4=�@�!;�lo�
�9yhS�J�e���Q�֥�Wa���M�3��S˔V�R�<=�#����<|-`��c①nh5�~�_��t�9�`I�,���)\1�y�U/C�G��E��_�B��/��U4�m��Jt��p���Q�à���t\�Tm����c�.��v��v�	&,�0b��z�M��O�/(�,�-J)�2��ڠ�'�q4��y�E�� ��� �, ��o�]��<=���us�1Z� ŀ2�/��'C�{�QBZ�����;}e�k��U�*w����S5�`��*#�Fa6O^��S�W��M*�4�-2����ɐ2T-�׏���$$�'&��ᘔ�|�tá���Yص^�C�K&����#'p�|�t C}n�~m���R���̫ƚ��|�������3��=�CAC���r�=�S�t��rI>���@\�*~�dI"��*s�
���7��3Tz}C��9VZ��7��C��d>U޼(p���� :b�F����}#��p�O}�ϵaݏ7��.nMN�� C;�<x;x>�yo��!��(MX�T��S������꡴�PuJ���T���,��j�,H����REy�)0�����j �U*��7�r�B�u;�A"�`96�MQ�#��
L�6��!��1A���t�e��\P�w.���d#�x-\fvIЦ�)@��ry�ŁviD�"�+]U�jMۑ�)��"J%���SC0onlB��mt��%�:����q_!a mǚ��0��$���*�^����b��ڊD[��m8���~��B��X�1�!�;/��@�N����y�ػ�D�ކ�آ�A?�/�ٵ��`��X$�],K|ʧ���W-��T�M��gB�T2y�b�N6���B ��!dV�C$��ͽGM+��0�
l[�9�i�W���}�9	�i0�ExdؚavaW�G��p��J�5]�w;H���L,kA����I��y�;�iP3����B/w%z��$s�\̘�O�~�V�l�M4���b�!���:�Y���&e�n[8O'�]u�ֱ Q�5��~����l#���W6���"�St/����E5t�J�Jd�(�c'w�b�i���W��'�~��/�F�9���n�h�'t9��ň�5Wo�y��χ���`�W���9�z�I�[׸��y�l(�a�M���@o]�	^{`>�c�>j�lh3�?�W3�H}R=S�˾�4�1�(��.���Q$7Xc���ȚEs53���%��}��-Pp�~]����xCt��@q���8ZA)�+;~���m��H��������`&�o�A-֊�4�n}r���H� �>eKFFeb@�Ľu�6[�Q4H��%����|�m}���xʅ�*���\��}�O����z{�J"eނ9����{�-��qw��|�<�M~(������i�>A���YM�섚�z]��}r��t�S�I�!�C'�:&�����Ԃ��n�c����`��!;��:�'v~���uN�&L�5��cH�ڮ-.�D����uR����<⧢��ī�g��4 	B�o9�M�< p�0g���r��",��>�4�NA��v͝��&�s.H�B+3��7?}�6?g�>l��fNAݦ�U���X6����MM	�힘3v"c���5����t�2�C�]��z
�pl���7�-���8�i�~������|�
6���D�頟�*��!�v}y�_�+��qT�q�H��Q�.�0�	�����~P�ׁ�(I��Ch���'�?i�	�Ӝ��iW�Y���{�6�;E�ڋ
S	5G|T���d~�X�����b�mb�L~E�oU���ܮ��do�F/�ffBb^���EVO{Q*��� 1I�,p�/�TGl�?*H�X�ۀ��&�����ıPy�S�C�-=�����~uN9�Kg"��qDucG��=CVC�O&H,u�zE$��f
�N�������O�p,ۛ��: J�=�. ʔ��, <�yJtC�,��W��8?+�t�3�T��O]������'N��Sҝ9o��y��1`veRb��.��/�175��k�g%���V��@�����RR}9�&�r¯_�ړ.rtK����|w��m��nϟ�u("���[��:��C%�7�P���v�J��3W��$nf��o��\���B�ě@Q�Uf�GK-������֟��`gਉ�0f�4��j0�7���2��T���M�Gry������d�=ܭI
��uk�¸��;�H#���1��5�3ڥ��i��m	s����/4]�� ���	?\|�.q�/'x�L�����Oc��'��ǥ��j�Ly�|Q��D�b	%�L��؀��"�X��$�H6��m겞|�2?M����#F�f��ܩ_X�^R,>j�l�`���+	��T�/_��rˏf��m�R��Ͽ߄���x����G��l�a�q�\�~��W���-Q�$�BPmd9�Ǟ��H�&����\�M9��Q��*�����S��e��n#I~�28�z��ԒI��Ѭ�w�YSK<?�&�t�*a)sw;�c���,.�j��б�>v�c��S�W �W�j�	B|_�Ħagj#���A� �a`�����T_��zDY��Kͨ�m�ICRyGP�1JW!��җ(q�|��'e�-\��Vz��þo����-���D�!~�,����Vޙ�pWG�'�=NA���}��
*Uv�x2��.��;��C���{f�\�8��ٵ��������Y5�-Ɩ�E����{�nIb죇���b��5��!Jv������8���
����O�\�1oAz�P��pi�=����_��>}���Uf�a�$���{���V��1	7n����A?���#rf���QZd�1�<��R� �p�xu'-�,�Ai(4Ⲑ���O��N�3u?�hԎ����ڢ�jп�i��o�]R��ՃK�q��Ar��:yL3�[����x9�l�JT�����{�Gd%_��=��t�%�m��PV�<|�P�R	:�]
4|
V��\s8҉G�qql)�b��]h��6��r%�h|�A�C���m!���D��]�Lt�e����]�^s7o�+Q^]�%�d�E�
`#��+�GΪ#I��=�Cᶲ~��Ab�Vъw��;?f�)��0n7j�t^W#�昋�8^����g4�/܊kZ�<%?5���k5�$ j�ZV��	[��uN��qt�ݕ��Mjf�%���qc�*c��M����W��DBX����-9��r!\\C�5�D�w'T\���32�֝{T�o�%��v�?c�R-�f�;N?�I�'z�V�M�v���A�V���a�"����Y6�V�zC��7 ��h)HӜ�c����.�ϐ��Mf]Qo�ƛ�+W(ъA[v������>cVG������N�2����J��O>I�!}/��S2H�E�/�3p�|!�HeӺ��",��fAS#t/��2�]��!¨�TB�[�e��m�<+Ge��C���慑�
!��o��[����$3� �hH����ġ�*\�����c�u�ByN���*�g'����wtց�a��*|	c*>�RX -_n��W�r�Rp�Ϥ�T�gim%r�΋�a��|,��Iu|��g�o�'�t�VU�"��:�ĴJ!��l�O!��cB��G��ܝ	A�b�������[0+���Y��muN�1CԌ���\J@�� �_F�r"�7���&\��Y��wM��j�T1�Ш�d�G��~(,�K��H�>��QW_�^�$&�S�7���fp�B�P�O���zk�0:�� �׿�gl��^��6�`W9���|^4��/r��.��z�ң����vI�`mz�,E����hj)C�nQK� Ǟ�OrG�n��w�Z�60`K'�����41���¡z�j��#�X��:��x�w���j\�ɿ��=M��Q:gTDB��%��&���~�_cA�y��9b4�CJF��6a��`����F�9T�ѱ�T������Q�%���⸉��<�X�ǲ��4��j�&��9<w\��t`c������d�N�R^@��S!�i�Ɲ��g�@M㍻�B��>(�p�2zS����6g�ӕ!��hё�^ȧ<G*�9[,,`�f�;��Y��	��5��r���R%�\���I'`�Cc�H�t�n�&�{D1��J�E�&��U8 �A����CN�B����ݼ�~��7��&U�����RN0��!���)��ǃ��և����p�a�C/1希
5�'���{��F@�2���?��?���{��������<��ۈ�޸!vU�'��l��aůcҒ��`��`��-_� t�õs}�o.��u�Sڙ�{&�e�g�ߧ8� 9F��9n$�ں�U)t��(�Y�?YT�hu�u U��:2�:�?������/Z����������{r��od������b����Ϲ5��+� �ug�_Xl0V�u�}2ӛJ��� �P!S��`
��Rg%y�=2ʞr<�:�����3&����� &��>��"U;x3����i/��#�Al1<�b�9��H��{��`a�� s5�tc��w�[��bq���کl�J4� ܠ+�;1&ZL�!���z>�-7�Õ�8��k��Mc�\����혙��X��5���Mg�*D�P݂����B�.�x�cV�P���I[�<��,�L�ϱI�8h_�x8t��Z��NZa�X�6�&?n^��t��E\3�l�a���BNrd�M梋�x¢��p�D�|r�|m��_ɇ#���F5׉��u��<j��v@;��;�+H�:�qb�'L��c:��j6|=�8e�
�=��{��cҳ���u��kb���A{ֆA5Ei8گtg�����׻:>t�t��NO�U��M�0^a�k �����^z�o��̩���YV���X�b�����ǎj��#�����Q�z�?޻���%��q�Z��j2X*oN~��J�S`�B'X�k�m�~I��w�J��LiC���W�`��F��L�]�x�`A�n�M�i,�8s��D�pM��L-0��._��M��H@fD�9���H	�٠���/ڇߺ(b�T/\�C�����%����%'d������І#���צ>����\1!�Q*|��;y���W�{ۗ@F�H�U@���9���E�����ƫf�4�	Й�T}��Cz�J�߲�]}�C��J�!/b���X&�E�
~.U�w�:�pޒ�X�,��DgF�񸩦��չ{^�S�<�i	�m���#�Gu� 7]��X|��uR-Y�!�=�?i����J4m蝓0Ea��� HE��_'���B|O�b쩵', ���;}�9r/ 3�F?{f�RB'�ib�:nۇn|ܩ���	�b�b����[����`�y���	U=NgX�4=��y�Y7�;�⋘�-�k��7^��B:n��I5Z �R��)F���A�63srȫ����3h=�E�+]ʾ�px/ �����������q0$ ���.�E���d^�	� �k�]2�i܂K�,)�ƝΌ69��ϸy������Od�BD,����N���S�OͰe[��-���H���.<�?��js^��0v����Nl��d�y�4�L~;H�e�I|� �?� ?��R|�Q�Or��Y���Ț���f)�V�ł]{75�"�K���e�w��ΐ=W�r�d���S,�Ok�����]�u���Ť�
ϥI�Sh!��������lY���u���aA�],�~��h��*�.�X��~�>H�|�{��㨭=��l��[q@��je�r	�.��T7�c�p��T������kF���
�T]U�Ǒ�N�T)f��*�?�����?0mBo�!�?ĉ}ރ�Y�����+y�N�>˽2�1R8{���I��}�S1i�����E�O{m٥�nN�MQڀ;�4h�}72�h����h����Ԕ0R�>u��߹P"XM��PfiրҾq~m���^�JJ�����c�Hdu=�O�j[/;t)�d�>���-�
��s����;,����ag�Ejȝ��<����h��ZO�ŭ�ₐq陠���y.ʋ�*��Hȅ���s*ڕ?�oV�|*}�6�����8�R��D1��q��F}��y1@9�g�W@�dۘ�P�yB)�5+�9ch~�Z��rE�K��@�.��;[�.?Mk�5��~��	 9ƭ��$���W�����`t�~����8Q���Rp�IqF=Wq��p���͵�c���L{[x����<|����{�^�����ʨXa�#L�d������8��{�(q�d|�ţ��ӗ��.���#�B��ˉ��ߩ���5��4��@�b��D�U.(��{�ԉD�P�7bl"�䌊[��i�v��8��i˦����>�e�lv��� f*=�%�S����Od���S������v���%��/�L�FIA}�UşI&/����d1��*����X���Y�@�U^����ZAC�-�����/2Q^��:b���� 䄹�@]�0J�;x@�A��3�G�
͢��'�;��Ȯ��jupiy;��嗹��������eb��M�F�	�e�߶v�<Y��Ʋalm����i&ڱv`���~�˕K�?��˛����ZB�b�˲�����½�|Ty�m��&��t��&,�陋
�n����_�K'�˅��LN�$���i�p�A�@�&���3�c�׎�$�(�a���p�p.{�q�nk2Pr�Y��i�����rl
8�cn���iX�8%$��5�oTo�i����̺`��T��;enJ�?YpY~�z��T�/xӐ�#F�;�_@����v+KHs��H��9�(60�1�1W���sn��7�L	�G�L$��E��LF����̡�j�����N���Y4/;��D*���|�0B��j�ŉ��P�rc�(��hH����������/�z'��H���֢�̿�~��eevn+�h�}	7���\QT2���V#��|x��w�d�,���]aH\j	��s��tBGi��n!F�cXI�ڽ�(��3���o��HG�ܢ�=��
��c��X ��q�gG7�0�s晻�����4�D�f�2��H�5AfS�x߽�F�{4�4ص��9��g��H��Ξ*���#�]W�(�q(*pB'���No���`�����-9���/6�z�"�7&�rXJW�ȓ�L)���<ՠ���IL29��pr�~I�w#�K�z��H#}��}��K�.wp���<s��s�>�ϞV�5hAP#�����CC�L���{X�:���Ṃ7��nu�^����X��z�'�D1/87X!a���3X%i����a'��Cl�.��nh� ��G{/+x�L��#*�NWꀽ�zbJ�g���S�Q���Z�_�Lh	�-i��1�ʧ3l�/E6'�	����{"�*m��E��GY���}6��հ���/)Y!v^�V�r� �	�zWJ w)�Qy'�g���򩒯j�v1�\2�>3��:p{�/b��k�(�iU�c��=����R������&��󉨩����3�
��"l����ډ���������|^��=/�ic���"�k-+b�g��.�+�X Ѥ$5��SV�@^�i��0x�AN����tstI(�Ĩ�ƣ� ����0�  ���ד��K��,a3���w�Y$�~��GS�&.g�bׄ[���ܮ-1��d����g'$�?��^�xo5U��{����mиR`A�����T]��0��8�����%�4w�a\,�64h����[3ڍ�T���^��P�GG��N��7-��ʡ�?�ꑉc.���*��D�p������pd*`b��Q���kNƕ&V��V�t
*�u�	8���פ��Q�
�.$a�t(}�t���;n���������s��fk���1҆uZ�)��RT/��$q�5M;�K��N2��ԱHN�v�x!����M����ǎ#mg�!b��Ro!O��tȿ�?$U���*��Z�UW2<&�6t�G�+=�R�D~����h"�a��[��0��D#�67G2���BpJ+��|�a������|˸�H��y#�K�����L<���WG\9�*:�e���q3��w��֑`S�
��\؜[TTO���<�c _�J�qp�g����˗O���z�"�PֱS-��Ӡ��;�pc_O-G��3�3��).�1�x2jכ�y�23ց^l�nѳ��w���Cd�7��ռ��˥#̾| �P�k�������HԆ����s�;|PTRZ����Z<7DD�zGKd毸���G58�%�vMOh<���2˙�-kJ�-U(_�{j���8����uSB�Z��0���Sb�}W�Em���g�c!nc���&������,#� ?8��R�������:�>��cc�4͕�yV��w��t��c�/.!�Ɗ�όK��O�r�P�f
�#ݘ�BV�[n
�2Y����̗ag���_�i��������ͬ��{`��_�BhX�+=(��n���pl��n1<2��4t��zY}}J�����4͓g���J�u��W򒚼�kZ���5ၶA�R1�wc�T>�_��#ȩ~y�^ی�����^2���Ѓ�T�e.,B���G�)����@`F�U�.�-�K��� ��bqPl�盻v{�v� ���tZQ�5�a޳��ԍ�|E��;�W�Q	<d�~܌i�wAiB�ۯ�U�����BH�ϝ��.�쵔8ǻ�(j�yf#x�-H
b�B.fC� JO� ���1��9Q2����J{�?#Q��Vl�O��	�O�M{�e�̧Atqz�c��-)����?�(�C�n�w��GO��a0����A��d��M}�FT{/05�ޘ !���ջ��Ho����g��hñ���NAL�A�3j�o�R��(�R#�G�F��N`�����9�0L��@K�D$�	P�E����8d����jM>"n|W�3�U�l�� a�9����܉{
�.��� �E������^�C����Y�m�q��?CƗ�i$��F�;d�R�A����1��+�*0�2��ü�]�O�أ;�?I(d!�|3xd��e<6���غ�4_/��3�緖VL��K	W�_:��Q��1�]���F��.E
z���ܨV@/j51��
��wK8��:!���U�-;�}�B���-/�B��U�<5W?7�.v�pn[Hp� ����V���a�+����+ǈ��T�V��R�=� V�.�4xHV�֯?��N,{�d���_��N�7�s��4�<��ͿÌ�I�����5�+=��V�y�F}Ǜ�$}W도�KB��Yr98u����!��QB��ڈut���1ZzTP"��dD3,���
W���|}@'��#���?��NKC	�6-g`�+R_���>����2��9�?��m���d��Nƭ��,U���Tg�ު�%Y+[�ô���γR]��M��u�eD�h4�lg�6š�
�}��L�(��(nѸ�(219�����R�9�u1��|�i'Bk|>��v�D�R(������wtY�z��[��p�e�|�qY�?�G�����!����+#�\��h¿�W�v�����t�CB�;����>Y����p���8C�)�@��c�����b��dw�V'��1�NM=�#G��g���W�	��*(7R�3�@�N2�g�9۾6L�ŴcF���]��\)�^����� '�WԞu�j���k�*��^T��.�>�(��w�I��=k+��=ľ����G~���.ݛ����Q�"M�V�d!~^ݝ%�w�&X���g����m��M��:�7)N�0I��$�2���x��-]H7��? ��QzDڎ�i�+I�hg)� ;�d���:�xt�~�q�QK�.�ǝ�yq�^��T�������M9C5H;��W��Sg�H�Қ�yY�ݱ���-ɫʓ�R��?BY��%�5�<}�CĘڧ��6�����2�݁�lx����S������f��1F��21g�L��F ��+�g���*<�PS�{/���Haz��/�e��/k��Om�<*�X�#�]�_�_u�/f'n��O�S�E7����r#I��e�:;'�h#U'��w�ƹe��8W�W�9`���� �t. �֝�=�	����4N�5ב�[�SVV�'k;o~"�K".�25�o�"�fZצ�T;me��{I0���~���:�b(b|u�B*������ia�ΐn7� ރ";���o�r븝���"��N�/K�HYd���5	`�V[HoJ��h��d�M�*�G�lȣ��{hIn%�}A����>���(�x;or��"H��	�b���k�.}xE,�lY�6�bJ��G-y����MgB��#⃢g`�%����D\&� �U	�w$���pUR�"�X΅�:�w�d-�&�l5ʦ��fKR]��c;��!x�(G՝�I8���cf��Cv���~F�d^��i�8��P���F%�3`����Hz6{����ӛ&3�wX��^���n�d-A�ξ��S�͐第Z�%���s$�CLLH�����v�&��][%#v�o�0ӥ1A��2�4H��� W$��F�Hkm|�?�(��#�as/쵕��̧�7~�� -�/s��%����B�kr��z=�2ң��B9�x��yQٕ͢�)#v}�И1;��hiZ��M�b��}b2��k(�3�2͞	F�"����N.-��6��/����6��Ļ�E*)�H���f"��9Y���ƺd\{�Z'���e6�y�·�oB�z�A'⢊��>yW2�b�o)� ۠T?����חW��n��܋q�Foř���0Gf�+bU�G��S0<�wνs\�#�]	C���h�(�S�	Q������ݰ$,ꦇh�Cs��f%%�~�ۻ�=���Q�|Y���$� �ث��{��ƪ{�S����V�5�`dŷ1�٧S��\�$+���d��N�-��*���-��{��ݧ�}�P�
��H���%�)�ac!NC��g�Λ�e��P�\-�̴[R�#)���1Ս�nu��q\4o~����k�
+�_��!�F=���!1�s���ӛݗ2|��b��o3iG�P3$";��6�9V�ƥ�D���w�@a��*���H�goj�3��ѼeU�t����I�co��跑�B���Y�v^sM0shQPb������s�ЍaA��������06(P���պ�byVAO�m��1��e�@0��ޛZjܤ��Q>ؿ��Ͻ��R�#��#�e+te��}� ��u:����9)���b��4o�VEw�G�cȞ�?A�����E���D(����a1�evV
}� 2k��\�l�,�{�� ��P���Dz����F�ţ���0__4S�j�La���ij��"~�cjm�(���a��"�����5��^�u�)o6��Q�6���A~[�.��i���G^�QSg�g��Z�'Ynѷ��vZ��3��"�X�7:DMfi��mhf���h�$����	��z?}����ؚ�L\����&ެ��O���WJDA~Mٳ��j�x�/�W�A-¿���gL ��n�|�z�[�{��Ύ
�%�RH�Oe��y�%���4M���� y��!�xyY�����<SX6�����h0�1��m>p��;��0�ޙׁ�Mq>�Z��H��}�?+�Y�Hbא!`<����4R��.�a�x �l�93:�ϖ���e1�n��5��-ʚ�O�&@���:��A���e������16���H^(.@ F�?{���%蕺���u/�K��#�#��{>|s��S]�o��A�+�k��`��4�6�OC��Z��AB2<���8l�@H��LI2���n�Y9���n�4<^I���٘���Ah}F�"�F�EŇ��8�tթmA��ڶ��=�0�ñ4N� i�pݨy�.���\�B,;~\SDY�����G���C����l���=�t&�}�U�!u�vA/ #L�G'�0�1��l?/6�G�����������})�1%��yB��]\����y�$ҁ���Ҳ b�r��P~�߷r��0���V^���L?Y�^R���PkNx|c��B�Ϯ@q�F0Ĝɍ.�m�뼔SIӍ�����aX:��C��^Ȋh1����4�h9���tx,3Uţk̔��]�׳�N4�N1�j쫴�F�B=Q����v�d�ׄ[�n���r�eH&Iy����|M�<Ñ�h�0�uo��woh������[��O �4�~����"Ylt{�U^�����l�F4��öu�R���K|�
)��$�z$+O|�{6�e���|��qk��)���τ�_�JS��|�y۾u��-(�nt�m���5h� ����C���|��q*���ّ$|�ngʟI�ȩy�g
F��
�h<��t3�3[��-�!�i��a&�
�>�7t�^aC�PU�����p�N�g(W��>.;:�.���'m	۬:��2�[��^aD��u��I��$�v�U��փ�uo�M���M��?o�ެ�g���eӍ��.w�3�ئ�/��X����u���k��S�/��T��-�B����jj HwNƽ�޲�0��i%�����~�e��2���ຣ[\ȥ���*�hd3�gA5���������Zl8uo�>lQP�y<�s��1~���Ӡ�C�C0���͑�)��{�+�CA�e$� ݦ\�΁�8�=D�������:Q��G��LYd7� ��kͷ�|µ�*��"�����q���zZ�H`�k��ȹ�y��O� ��9й�w�ߘ�ӒL%'	ĉ����o���y<��w�2\�z�)�
�E,r���Z"SV��֫����}M�Y�h A�	�ʳ6W0���@s��#�(�f�|�����2օ\ʞ�ܵ𣂎���D��*3�V�Є��V?�㘁0A��)�����s����["~��P��Z�#;M|*�Ǹ�k��c�,V��*�3G�Yq"ܑ�� ��e]�Ӝ�g/��)�4 �±#��YT������h:��k��Aq�W��g�O��� F�",�|�a�p�o�^sU�-��_���s�ZlV>��M7�����'�h�L4��ZC_�.u�@�=-�;6����!&�9���]
��a���`�T4ܣȍ��h".�\����ʝ�ڒ��2����]E@�y�	�6�i:�ؿ�y�sW&;��@=�{#!g�q�
2Ç_�'�8_g[�fْ(�Q:;��{��,P
��4.%��n.��}��u��@��@��1�|��G��N?_��E2L+HS��~�c$P�u�����V�/E��8�{��O�qD3���ڻC{���o��kg�]�W36`�����1�:o[�b��ٮk�S\��X\�����Zw��b&�Ѓ������X���a+%G͞�_:�I0��튖~����P���/�i�^�/�̬\���z��H(4]	�F�G'WV�!0?cI&Es�`�%�E!@
���䰖��]Lw�s����?[��X�$c��.pWi��Ī����׹�� �Ǖ7�����2h65���Fj٧�_�^�3�mW���BB$§/��l?���n��2��L\�j��OİO� <�'+�B����%*"x�[9�L��q����H~�7�g�]j�M��w ��F|Uﲩ��x`h���ٵܢ�[�o<d���Y��P%G�EZd��T�n�����P��g����;���E�5L"Hqw���R?+���v6�#�&���5PCq?� �)>E��P��3t"윀��u�L�0ȭ۷�H �_�/iw�?d%+�����[M8d��+)"?Wh 6S���;{���L3`��|�N�u1�v�H��b��LL��O���j��b90�N}\+�ŧ
|+�� ��ζ|���g
['�U�Pb��(�M���FY�ŀ����䁺5Ә�z���a�/nj�����ʿ������n���y��
>�Ͽ,�����'Tn��i%��=+�^b��z휠(���v�+���tHN��m���r��5��"��Ж?�-:�B
<��9�1;Y�[3ϒV��ͺ��%�(@K�s"d�V��l���w������t�'�/@�6y'o[sg�7I|���(aM"K�je`Rv��F��K�����zOdD�c=nU\���W+���/]R�U%?�9�6�b�c�,q%��@���.���ʦ=����K"c��V���8;_Ap�iPd⾑�.L �kHȕr۪Ծl9Gᷧ{?*|*SXA����h����!��=��.�
UЏ�;��V�����ZIq [�!qU����M�q7�#�~T�?�(=2*u�Z�������ې�w�uZ5oy�&��ZTh�tB
>D����u�p�vF�n8Z��<(��fU4"=�?#�ꉏÞ�v��i%�?��"~����9�Z��f�����#E��k=�j/�}<��Ў]9Bw��`�y��k�z��H"�!%����<�[�H�P����B���o�O�[_��s)�;���G.�#����}�ה�����rd�լ���_N,8��s#ڝ'
�}���֐d�kh@}�X(_ږE3�z� �TY!Q٫��iٵ�����D���N'�[9����Z�1�� \!����|07�s�����_�ı��{��@��"��g���`Rt��X�~۔q�����(��T����S���冶ƕ�~'=ʞ����^�w^�(D"����Q��3�a"$�E�t.����(x�&��g掂 �W�GN/�"��o���� ⿋bi3�*�ͮ C�`�n�����O �~��-pty��1@�	�J3�i�[!�/�C#�__nD�A�)�����a ��{���V�����rBp��u�Dm��_�-����,���)�d�Bc�Y������V�y>��qY�r2$ox�u-�U���v�'����2�L\5-�]����f$x���5�qd�i���)�HL�yf���3�qF�H|���mH9f��j��<gU�L��6���he���x�E�˗ܖ�d>M�E�a�l�a4S�)��W
�hX��U��-�]��>��Y+S�1WVT�z܇>HV��N&%\.�3Y�|���%D����@�tgN(.`Yt{�I���h��W�-Ga���m���=W�~ 2�&iKx��Μσ|v��PR����G4\b�GţBkw�@�l �
�)2	+�J���(��
���,ޤLt!�4�z�d.d��j0�n��+�~-@����X0TH(�$:��#�#��'�gU��Q�tr����kr�%��<	h`�C�ŏ�Z��_�X��7d����(��,�]��u�dl׏��ӫDz��ǂ[� f���qI�E�C���5OJ|����tZ����n����i�A�B��а��V.ӳ�3rE9���U<��1���M	}@���<2/��L��l��&���G�>�Kհ��j�n�L�ߴm*?���;�t:{RU:�Q0;�M��U�����(�I6޶��G�ƮG�
��Uuf(/��pA�gG"����ï�5Vh��S�ۅ����ء�����Q�‘Rs��L�=��wq��N)�70X�DL�"Y̓F[��W��6 Y�p��y��ꐬ��?͜�N��,�|�|��Z�˭It�Jq���F0x��kSM߾���>����,e��K;� ����J	\	�R�lh�x�@2Li�mQ\��ț@��S�!RXK���!�δ�?��Nۓ��t�C��7G�B9�T��A�1�M��BqN��nX6Q�`��7��rVY]8���Ϣ^ѧ2K��{��]�'�t���/������KߠN��em�%8�p��{����퇙���7{O@8�4'���L�A���\S���Y�־�CC]�P�ߵ��4h&B�3e�"�,S?��2II�����[C�u�����мmBBbĨ���ZK=Au��ٺ���&N~���"V�?\��wM�����68�h�IH�F%G��Y�<|!�)�Æg����$e�w�0[��l�(���
��K��
��¸A������N ��k)����x3�ɲ�D=r&y�s���:��'r
�	\�A�^��Mƻ�{��K�"5-�t�nu�ƎJ~^<�?�&�����[�<���`�%pA�w>^���Z*� ;��1\!-�aW�X��C���=5�)ANe�aI(�"�T�Rnq��q�%o�|u�UJ�"����K��- �L��F��f��<�B�Բ���%^�Y�9mi,o��3m@)� �u�#���9c���pѫ:J���!ԝ�"'n�,fnj��A�^�7��]�󮑅��	����2�y���0����P�J�[���&RZ�"��n_�U��k��߉^\�ӹ�1�i���=,y�7X�e��D�u���P�j�+=�!�_�8�H�n�3/�����h.:����x����-��J	א�k��2R�5A0����cl��K��@�M���y��c?`�k�^X���
�%��Ɵn���i�m�h��R���C�$k1�X�����p�������ee�k�}D�ֶA7I��v��9{���>WCuSh��P:=
�����]ஆI(��n���|¸\�^�����O���+�%>��K&��0/�����0š�T��b�\��ة����/��o0����S���!���=��{f����/����˞��J? �o�ƨ3~N��Je��M�rQN�d�D-�I�ߜ:�ޑf1�_���-���b��\Cа-O��N�2�9o�bJ�B5̧�8U0U��,>
6��~/�l���	�"�2T�5Wv�^kM�`�|GM	��P�Z�g��oZ+�ܝ%�. ��(�\���
��mR��r?�s��;8���ࢨ����U���a��a��F�B7�m뿏�In���6�q�<U���&Z2�l��|7X��),йj�cO�ZjJfp'��r���\F��&����o����##|�D�\����B��1ˡ`��@e�ow�5���*��9w�fAL��yp�C�Z���o�S;�����V�{e�Ws���>�Q2'uO'��ŀ|���i���@eI�%�b����cl�X�xy��f����F?��k��zy�d����k����Of��r��%P-���q�v;�ӊ%��O�&{���n�Ja]����Z����l0�M;�I���I�GH��.=��#�8������pUЍ�sd��~7ңИ�]G�t7���ib���`~��	O�2N���|6]�5��[a��{_M�A��uo?����9=:��g}��W��ז�Ot�j����5���aBcܶ��~Dڳ5a9˗O�Ey���tU�G��o�"*��1�&�^��.�ú�`h.�&�S�m����_��5dzxN1��Gֵ�m�/�Q���v�=\�@���Y	'�B��j-�.���DA�Kq�	u���P���7�Ů�e�J��D>���S'��0� 6t��o[�8G��;8�ô�xn+��6Pm\
����j����hۍO�#G�-y���	=���K��>�H�n�=�m���$ύm��k7�����D�g�*�=�\��t�Sw��yE�0Ͽ��bџ��YJ%�┒k.�і�QW���v�1瓮��_��#F��I�������0/OR�4H��;as�]%�ū��";�h;?�7�1�?ۍSuޭ|V�V$`N<������f����Y]����y��[�Q&�������t!L�T1ߡWC��hK�G�_�2����
ϟ��x����=�3�cA-^F�����Tթ��uҔt}~��(� �l(��u��Ⱦ)�z^}��Fj�:L�NL5g5JC��a������N��]HRd�/u��<]�_�ۢn0�1?�羶3azvq�WM[4�=���q��t"�=��2"�f�s�!��9��SC7�����Y�u�!�ًi������$J�]�z0L|�ϰ�d����U�b�C���������]Im�n��\�7��֝�BU�������6��-`�Qѫ
\�m����E���C[�w`5'>K٥\��W�@���Z���@�����UmvS/DB	.�E!"��Fw�$�a�Z��+�-�Y|���
��^�MX-���H�%�J<e���W7���ZSS�^��D4��/�1�</}'t	��l&�������������a��Eid�~:,AL� հ���/F�wY-.vں�p���A�GnK���38�|@=�@ư}2~���w��.2�ךz��Q3���JD�B��e�d��"Z�T�+)�`�9��A��U�ٴ0��w��Ǘ3�seI�C�M��m�顑������]``�������^�N�m�`l-8�n�ĉ߈F���l=@��:S|Cߤ�Ŵӊ�!����2%|h/��6đL��/�|� ��*����^�
��M3�-�&{m|�d ���>H���6)^�B��O���b��C����7rϜ�c�M��*�m�(���\"��50.@��� `�}�U��7�]�� ��`���	�(!�5��A��� <�n�4���5���U/e��eZr��cn.��#�洺GwW��V／�U��	N[~���EI��uZ����z�tL��7��O�~&G�]��{���&y�R��X>q}��[s�F�@#r�*Gب��;���|�*�U%ws��/��L�����c�Ñ¤tXyk&E
Y o@�B��L��c&[�ͨT��l<�?@�{��-SbO]p9�ñS>���"+���v�Q萶�WG��h���G�r��;��u/ޞL��L�5k+���4����'��)�	��ܙhy��'t�I��7�A�rf_�f�6�xIqB���:^A��T��Zf$��P�ym�&=W�
�����zɡ�tV_]��b��H����]�N[�< �v߿9�4åS�rބ�����U�Vm�s- ~
ׅ\>�F�k��7��%�����S��_���8�.T4��:��QoUͦ���|�ϑlh�j�}�����G��8�|Q�,."��8��j[��IV�&{&��T#����d	�[_�%�H>����k����Z.�z��J����el�'��I�%�cɢ�W6^�{��� y�z�3*G�P������6�i���}& |ґ���C8����'F2-��iɬr��bC�)x��C;�%� �xs����9��a�$�l/$H�v_4��<-£�u �{w�@8G�8ى��ՙ���ɍ.O�G�QD}�q*,T�v����=�ʁ�ܑi��ȁ��Y�a�7�zD��=|,ƿ���B�D�ݽ��HNL^gh)Ȭ7;�Z*�;V�<�x��I�3��6��ư}M�q���SW�X*���aA�Y�U����7տ%U��Q�m��/�!�čk�kKazӆͦ6���A���Xl�����!j  ������m�o�ҥ���R�3T��FY�æJO��?y�VY��rj�dG�i�,?/b�H�yF%���ح�o9��p��4rdd�?`��u�i�5Gd��ġZ��!�w;B�dt�Ff��4{ӝb@Q/y����CC��S�9�$b
?Pm�#Q��{]1p�S�4�ִ ���o���q��5�'��Q��nR�d�k=؍��0J��m=��O��>(��.�n`�X�L����Z��?K3�Gw{��w�h�d��Y�<P�V�e�M��i|k��Q��k��!�XC�W2�h�"��B��3;l���Aڤrҹ
=�U0���h�3�hQU�'��7d�Ȑ�L���Ա��I�)�W�%�h���NV�侞$"���۬s�D�N��T����n���n	�,��/$�id�x�/)��'�Ƀ@9�ʣ@G%���O�SL�����_��R�������HI.+;g�>��W���WQ�@t��#�T/�6�w(�!�2)�(+�Ƨ}5*�
w؈4_�Ln�?Y�z�܎�VF�}C�""�+�[��C�A�=fh��E��-GP���R�j�F��Dl�cW�����S�Y'^���G`����$[Ǧ�������e�t:d��"G��Db���Te�S�_�Q�i�ĽT�&��y�]��:%TP�D��An��Yͤr�Oc�Հ�5�E�oXO�1����];�6[�#� ���i�8�}�'0�����L���7H��� N��Cf�a�[�K���U��dEZ���d�����vt����"�(�|�W���TV�00YҮbL��:�#��^�F*1�w:��--�J�U�Āx�kGIbje�$�R$�L�'�n�>d��o��'����(O'2��+�r߭���>!]9������?�
���.\�Nó��ګld.��:������h���1��q*�g�Z@��qGc�� �iU�n/"waE"��VV'��ɾ��0��2!apèP��L-�p�n⊋��1]��@�wuR�sMu�{���6��
��!�v062H۱�5��ۢ���iq�ۗ����!?�������á�+������#0y�R@���ו�=�ٷ����\���K�����T�s���B�y��Z���Z��@�Y����O��J����r���u��`GAp���*�Tc�����5Nm1��L���Y��D/��zAbqK�9Ժ�f[��U?�	�ӏ�9�>d2���`7��nE��O�'/m������4��W�Ҍc�S��l���q�,�&�%ݱV!'�����g���1�w/�-\ �M���]W�n7F��'��}|2r*9���<Q8�%�m{�s�����?R�H�1��F-��j��Óu��.�8u��,�Du�M��mw�<~Ӯv=�NȚ�z7���wő�����;Xx �؜m� �-O�[Z�k����Ŗ�dr�X!)Z���:>{0�D�1���oa�w��G&�#�j+�f��zx{<�Wqc���PW=�=	w�.j%������kw�g.�I� �͆;�^��Jh_:��{&:�)-&T�3�Bǟ�+\H��q��%7�3�zJm/CrV
}��[#�;~0�B��$�y�!��hx|�t�5۴Og�V�ĥ+��
�+�|q,��k���녖U�X��ۆ���BÌ�ن��=���[q��^�P0tb�߶B�9t��lt�Ȏ����i���IP!��.t7ٟ�BA�i�����Yy��g 1+���˙������g0�He�Ϗ�gc�$�֌2l�-L��Y~�/�N��s����"�cݼ(��7�S��m|���$��cϛOv�粰\�(��J���Ix����8Ht�tP�i��tU�$]��M˭4�LEK'�)��?�*=	�N=-fQ�?o��G�]z -�`t���&p_���=W���!�0u�O����~]t~���];������' m���\��x	�V����/x�*�!��$�^z�J�:�f?B��H&t�g4�����Z���K���ث�X���df�d{W�ׅ0�\�����z��.��dl\�{C�]/���D�TLR^�L0==��ԔpV�"築&#m��y�����;�[Da�\O�KK���>��#C�ʌ��9�Н���nHt��auY����T%`��-k`��y�bƜ��� ��&�!�<��AD���@N��5ۨgp4=Eٔ����i:�eP8�|��s�^�6�y[��.qR~򂧧ߌ����#��sy�����J_���	(=�sz�>��HV�u���f���,��^ٲ"�M?��\	�(��W���M��v�ݥ�6�ᢧ܆����Xs]&��i�����ʈ�U�ib�rb��qK�&���銮ʮgy��_���!W;������S�/ޞLq2����U;d3/ّmA-��2��`	�b^qOo��}��O�k7���"FIn�
ۢ
a�i�|$��hP�7��l0�5�Y[�ڃ\H!a�-?�8?�먏h��D���Uq�(�)���`�3���d�&��u��M���Ȗw��W�W�gڨi%3P�� 4����_�7��a[���]�8�CDG���o5��f�Q[z?Y����\�2�2��`>`FZ�z�?�Y[�dd4ٴ�?nE��ôZN;u���_>M�$����c�F���]�bó�Ǯ�OQ��#�_{GM�ᶱ�A�Ş+N
��G�+~�sCNev1�J�g\�~ <�_9�9�yl4N��-�P{��Wd���SpT�s{�^IY�<l�¬ۗ�ײ*2�i�5,�጑,���r��|�(�ϩ�#+�����OrTO"������3�C{�du m{Ah3r�o_(Z+�����ԊzwN�a^N���zrHy
�,+��x�ו��3�b/!'+(��2�,�%��e�،pS��jN��A=p��f���ϧ��ka�SJ#$r�Ŋ�-���y����k�@w�2�d� ��X��@':�S��!��֏8����!��k0���N�����K#���(/�Ց���{��ag�jǝd蕰Y�����Y�T;r������0�U��/96�'�_)�x��q\�{��Og+"?'$l��	e��)in�J�%�]�Pd}�.E�f�H褅� '�Y0���/��u��Nbo�)%�����%['\a�2�Y�"K�3VF���P�s���-$:���	����{����J±���O�Tk<}pm'ȸ!�qf ����p�UH�mǴ3QWW�R������C�"l���&�`��'A�ֈ�A�hn78������:[wPFS�u���nrN��Wu!���<�xN�J�1Eg4z�ڕc[ |S�^yl�6�n/}�ZUt�D����=�ocd�����^�/9;Y�xW��C4-?���b�Z���� ���t��>˞h� +kEߡ�Ӥ!sNTӀ��
�¶)��&����m~&�6��jQ����Y���ʄu�[Ix2�%f��Ky)^
��W[V����[�Ü&��l��;VO$�}�Y�bv� �&��C�4�����7���h�L�/��K	�V2\����Ga�IH�̻�ƥ_�y h����!�L�~Vc� 'Xj H���x�>Z����\g=�[�}����b��r�s0M�y��t��q�
5-�K1гA����͌2�8G��� �7�vX����Q�����.��(=Jr�"V����=�E�M����`K��d/��ւA����;H��A��G6�����f���%�^��G��`��{�6*	�y��nv�CWő�(	lg�J�ʱ6g��=���&ڱ28����ԯ�Y�.t'#����\��ּS�(^���?���I�k���Q�T�R���,R2�O�,����fPB���uapH}b�7�y����D!wC�W��`�*]i�Ì���w��#����V��T�5H�\$d5U�����v��L� BZ���;��Ob�2%ńPYqEi����sҫ����4h(<3��&�={L�����~gʧ�s$c,�c�skɢ�9z�k|zx���]܍L��m�%�1T�o'F^���s2�Y�72u����b��q	^��~��Ĭ��O�s��C�Q��_�-j�!���t̿|JW�=���jT�5�MI�w�{�[��ݖ-l������|�SD}��t%f�͇rI��zVtt���g{S�P���(hp�t�v���'�Y��`r��H�U�I���p!j-l��myh3*u�Fz�f;
N�1��<ρI�Y������<��Tu��=�ݕ��ak�r$ӥΎ�OO�Oh��2M{��m�Ū�M~���NH2������kK������ύ����2�� h&Ҏ��~��	�G��C}�R���������Oa�6ɉ���:����`��� \�K�Ek�u/�BϱoeY܅b�1�do����kF�n��a���q���c� ���P[O�gJlb�!�����=|(�o�{Ҵ��l�aZ�.f8�7ZV33�I�q��ߌ�@�u)����ɸ����aK����
m��eD�PY@��7jS��v�iv0��ȬI�{��PH1���m�т�Zy�fШ��mx�^PF��u�F�!����|)�����ރ?�}�a���!(���/KzF5)4Fu�	ڇ.�L=066\e���kyR��U�h 4^�CD�'P�*K���u�l|���]k��]~1Ԁa5~�T��W,v�-�W���[�	����	���̤��_7��]9�>Vl�=MP���_�.���e�U��?o����f�*_$����9�׮(/nxF@a�m7͵��~"^�E�D��z:�3�xƺ�@�/��٪D@ҐD�y���Dw������v���P��X�iI
��
U�wh��Jc�b�=h�RlS��y�t�0�~�D�0��&vng���.��х��|�t�¸�?[�x��L�ݻ�('b��k�'uVvgAv�&<�����{�r��d7���#^2�fEټ�B�9��Q��Qz/^���qV��v�۷��5�bK}��*��-$6�N�\�B�W�����?*.��oѕ,��<���VV�M|l�����:#��/!��"�ƻ:��u'0�Q�\�;S E*�+�l�-\�uS�g��2[���,rHj_���X����t�[�w�O�d�Lj·^O����������T�)�M�/�����(|�2��?���d��i��}9�R�2�8E8^e���i�r˾�KU�類r����y�G�-A&�7n%t��n�la��d��5"�K��!i��v`�n��s��v ��=^^�j���dԕ�[����Ruc���`X�����s�	��*pc�ӛu%G.V��b�|7h����J8���~�3��E�0q��׹XEr����=�����ɏ
8F�;��kS@*����2���Z���L�o��'2L�����g�>�Ҝ-�x/����:q�P�N)�o(��Wf��%�w4|�׏����8�I�W{�sն�����Y(n�Ȁ��C�7VǴ.���ˬ��W�W0�(��)�U!��XW�/��Lf�����kAޥ��j-�_����:҂d���������.Eq'k�X7��*���9�F��;��f5o�:�� �m9�nM��2b+l�����f7t��cT�/O_�$}O��$��Kp�U{	j=�s�.M]�OXc�we�,XA$M5�uLZM��\��ә�(d�)y=�.,V��xN�Ϟ
� 茶��,�~��c~���V/'J�-OH'���#���߄��+��҆7�#\�J6�ك~L@_Y�����M%o�۳�.a����
�R�q�lo��\� ���\F�Pګ\�u�2��g"&<�Q�i�m�I��E
ֿL�t��V����[M56J��x���ǡ��r@���K������ZL�(�w|�H�k`�ƴN�n�v` �񭊱�����\(����s$���%�M��s������ kM�;�X��; e0��	q��B��v����HP2H>G����٧��bkB4��qq3s� @����m��\ �=��e���|�	�(��*� w�8��"�\Ϧ��C���#M��`æ9'NɃ=AB}��#�,�?�k�@5PY`�DLH���b��[R�J�ٚ���X����Yrz��D\�-6a/�n9���亃?n��\��1��_�(���KGL�G�G�~pjp6����� ��[��DE���=��Ed��3���΁�=�P�ī5g#V���GS���+�s.#�{��6qɮ��&]��b.<d,�R9�Q�T�n�ߝ9�Y�i�u�/�IU>Y��Q�]p�n۾�ҹ����%fJ�x�	z�lfz��/a`�r���	�T"霼�f#��	�?:���0Vn�O+o�4��*��b9+�u�fFw!ٸP:
Ja���N��J�h&8n�I�~�9P
.��QtMz�Y��U���;���e�B�OE���w�Sס�Clko7�O�E~\I�V��a ��6�/�=H�}w��65uF��,��`��l�߮��q����ؿ�;�T%>_H�Bc���<�L!S�v��u�Z:ؐŕ�BhfE������h#\�A8�C���I9�?�O�P	��yH�ȑu�	��$�r:g�s�����O����%Uu�Y_���$��W��A��U���k���cE�A�m�f�b�Š)� l�X�֨�ǫ�dtG�l��B���ڃel�FA|��>Fs�x�P��jq��O��ȯJ�����|��W5�\��u���it�	7�c'3 X-ݘ���X���� [-�oej ���h;�Q-T��wc:g�l���}���%�G�N>p�v��p�~?gm�"qmQ�T��@�]�� ߠ�!=�M`��J@�f�V
,,�-��iB3Ńbns�䎾�~]�դ$���o(eʄ�\ M������&N�Q*�cB�_��,���D��h �f��%�l{�S�Y�A?0�G�;)>Դ�W�veC8�e%(����o���� zm�"V�T�	�=���~�K��ͤ0��|��ͅ�������<4d�[^�n/免�KD��)�Y =T�6P;��#��Q�T�D��x?�I#'��COd��Lo�����@�H=����R`�~	I'����=���"����B#��������\�QK~�s��*1����gS%]�6(^���c��8xsVUoNJ	ua9�)�@�~ �bA�	}n�d�Fh��R�5R�� +��K��.�B�pʲ�B��4cm�m��G0<��Pl�t������!�6�e2Xw3��)��E>j}�������n:�x 3G*ʌ���]#n$Wf<�s%��A�O��9u�lb	������j��y�����Nӵ�e���TI�od���ؑ���Rk���%�WAr�h>"׮�o�b?�Z�\T��ǩV�A�e�z
��,슸r��d��UWey�+�:�B���rq�׊2���U�rIɚ3A&���af+l!>ߍc���eP��+�r}n�{V�5U��W����*�bYBr�-<؟*+�'|s�;˴J�\��ņ������lb~�9� ���$G8s<��T�����q�6�Q�/��mZ;4���m�a{���4W��C��}ݒ"N��.�!&�����n�f�Y��n�`+��B�գK�L�C�)i�V���~�_xA�J��r_��z�\,Ư]��=V���%B�԰��S �>e$�0�e�&!��9d�+��fz��Cn[M��tU�@�����>���7�,%y����}FC3�/)�{Ɂ}�dUS��]K	d��&������|�tѭ����L�L�i8I`ȴYeU5��:��KzqT�*�*��'+�	V2p��K5����bN��:��JG#lj��7�����^��K�aH��%yX!� ��P�f�D�F�%�O�"[K�$�.3A�ڰ�Q\���Y�!ҭ�$(��	��$�rXuD�ȯ�?�Cx�?�W���0}h/��p����t�ZQ���*3y�E_��ݔ�����u^	{P�o���+�~���&��C�s���o�[E�$�r�w����t��_aۥ)N���!s���[L�u}T�7Ni��U%��O��W��)�� ���qUK�aֻ�3a�wp�YzH x�P�7�w����l���D�t�b��l��E5m�7d'�]��B���m��\��)P0߇��i�+�j!�P�+K��9�����%tJ��~��*q����y��7�Z�Hj.�CH
�EE��	ļ� �pujIs*�$!vnϞ!��9-�l�j�#�Wl�3|�oȈ�R���iV���f�o�o�˪�vP�e�'}��-"(��r�zI�`��&hwu�*y�8/�TQ;R�?��$��G.���-���
�kթ���u%�1��%��Qj"\7s4^Wj�Q=l�j(�
��!eg��+Р�u�
>��^ �>��?���S�:����_��_t�]K�U���,&�Fd�',1K���r&�ٞ��g]+�*{Z}���Ā� ;c�-D��Iv7���6�Ɋ ��}1��A\��@
�y�W�j��4'���\VLܼy��~LX$V�A�1QR�`�q�y�~)&�Y���cg�L�!W�ؒw�I��7j�
���%a`��ޙ8�I�B�����n��f�t1���>�A�M�i���{oÇ���Ϡ���@g���u�͉��i�,.�����L�TC��s�5�C���������E��]�=����wPоA�A�O�z�O��L+�HVu�^�x��!E8����j���ժ��ǣ!fk�I��g��������WNL���Wr�%8W�����-pss�|�|+��/��NڦA��J7�#*�4�����"4i������#�S����t&���.�&��D���\���5�>"j�ˣ���n���UAc/�&3oR�*���z��9�(&��"1�O^4���e�����Q�b����-��?�n�H����ҲX/!9���Q^��٥|j��\I؋ޫ����svuѲ�J�O@N�-r��s+�Nj��cE&������/���t�����ӷ�UcL���ݎ}8�kR
��/`"*@��(���ЙN����=#z�.��{���	g�J��m/?�m�@m����H$��c7#�Ϛ�3K��w�Wt�A��y`������\l$.x���J*!��l�?�%�
v�;9�#�Ⱦ�f�dW�o&="�Jd��$z���� o����;PƼj�
���xw�
�T�l�mS���m8Ʀ�(M������2��/{�/Rf�$�)x�Ҕ�1���m�?�.�M����{ܸ%���Ş9��O, �jģ �^!��زG.�Q&`��I�;���r`����|,�z���M+<9Rk�{���N����+�
Pڏ���α��a���LR��9���Ӟ	�JU�TT�X�(��}��#4����eȸo��n�YS���?pj�|XkI1e;�l�}�91�(P	�qJ��I�w��&�����~ �|��eDH,�~m�5�T��`|$)���Z��B������m�ʇy�(,��7z�>?Cޮ8K����v��/U逭߮��9M�i�r�L����U��nF�O0���!*��/=1Ԝ��GIIB(ݾ�>���S�`R�R`���Z�5�A����8��#�������}��2T�^�Qm&��21�6T������q?��,�M$�==�X�*���F/H���Q:���l>U�v��Y��,�>���&�_�Q��Q�snf�K2���44��a�F��٢��pXD{�Xn��B�nc$�6��o�ωC�5yu��������]��O�Ŀ�?�)������K\��Vs��t�L�7�ޗ)x���@"���˼a��"/��:�E2K.3�y�r:����"�J̲��sp��ZS7�"��W��yl؎9��6����-S��r!��%$ew����_�%��6+�)"�'Ƅ����]�:�Pi�@>^�cd���/[y��[�w����bS�G�z9j�N������[��Q��!�-;ja�/3�}�%��It���N��:����n/nLU{��Dp;X�V��H�V��٧�bk���z��\"5��5�9��
z�q�Sڭ�+��������	��vȬїc5o��
�`{Z��Y���Z��f�iaMF�*84~I#� pI��Ҹ�L]n�A�$���Y���C����S�+�B�L�g�U���Y�V~�'����O�_�O������H�yӽ]�/��^�4�$���4/):<���\���Ԅ��m�t�E�r=��)g���/���
�?s-)�-k&������2�iks "���.�5�$x#P��mh��c�g|J�8X�}}儌_i�w<Rbz���]o������Ջg1���<��*��Y|3���5Ei:~��/)w�x�>7�'�EvȀ���N5�V��|�h��A��d�U���/��-W�j��a�
Rc+���N��)�\���L�zv�R�F�Aן�TE,$-]C����d�R�!X2��PM��1���2�_ �S\�<�j� �Q���N��3��`9���ڲ����W�TTፖWw:�[%�5u0�a�`䤢����p��
v�*���f�{\1�	zJ�N�v�CH��x�eR!�����P)�(����K�׼׵�֞L�0�:]�I �"ޱ3ZQ����""�7(S���y��ʝ\���m\=:����iB��RJ�m�������|4�Mbl��Z����O����T�ί�����k�h�W՞ ;��)�3@�d��G�м�`m���ko�`4�TpmX���ެ��Y�r�M�&���#I��]�h-���G$�>���½���.�6�1���@!c���F�A��1�}��b�&��R�p�!�N�vG��V�'�<2M��)Z��%�մ��!�Fx���ȴě��G�U��r�F)�T�P{�`��K[8��V1'���duMg~%�l�'T ��7�dY��)"	�� ��8�Q��+��Vtt��m���8e��,X��;��Nmp�l�m є�1���A�b!V̬n���0@�� ~�{�^���0�A��?I&�/�-Hqt�R^��I�b��v��.-�@0&�V-�Z��]�qQK��i����~&�P
�����#�O�_�ȗD��]h1%���眚�uU=;[����-���n$2V�9�p��yX1υ��Z=6'�H|e�3��	/����w��G�߳ړ�W$`?u�D�Fn}�0�C�ƌ&����;�{֎�v�'�]���3`�b�6�8�(�  ��r�PM��p��S�a����T��[�%�^H��P�'�Ɂ�#���y�*��PW1�`$m�l��D�{凰�k4�lw�OS�xS�[Gɟ_��{�Zz(#���m�%	q��Y��O�����iB��X��hာ�� |�J�F��9Rc����	�F^���_nN6v�[4Nzq=�~��|��)�\Ob�'�%6��󠐵�XH���|�=Y0�:N@���M5��$�<�wWp1���Hk���U���ˍ>��K]�N&���k8�p�D��٥+���~��
�F|k�ã"lW"6<P�}�w!�}$֏=�*,y'Rq�e�C{�a��G�����������k
e�Į7��fN�����F��a��Vn�9W�`]J,����> ����B�\��w2֫R� ��}�S�KS��8���T�'��:�MI~(ZܔY�?ػZ�
6�yäfR��#!ݜ�`�ދ�J������6��T�
68�Ҋz�	%��'���Մ�18.~&�:���)���ҺI��
@]�=�Z�@��GhB~�.P5ňo��n �˽����@�7ͬ��^�i�Q��p���}2�YV4F0SA���*��.Drk��'V�W�t}���䳰-��/�@�1�4���Ki�(=�7� ��i[�#�,�W�p�o�Br�A�޳��M?A���,�tK��k3hOd���i��\�c��U`�z]��x�������;ޔ[�(��/`��P��B�E��x�VW��O�Q�s�x�ڭ��O03sM{�SF);�	�I!T����;���]�FF;��W������<�D$8jZ5���Y�So��3�H��o+�x�+�ʩ��
�B�g���ݲ34;_x�-;���
yro��.�%؁��1Y�|��p,,�n$��t`�
K�X��$����B�9CT����p��p�g�>�9w�����^M�m��h'��+�܋���!��@CY3k�tp�.x�顕tU~��'82q@��͟�R���u�E�J����h�eh���ϩ2ve&�Ѵ��-C)r��=ڌ�h��}DȀD�;���WB�?�͵;��&�?J�94�I�.L�r}J��>�`cz$CW4CI���<��Es�MKΦw�i���ݐ��%� `�8
� ��:�Z�K��]#}�Nu�Շ
_qB�Lޤ��>凈"zb�[����1<���V���<�t�t�nٱ�	Р�Ꞷ�d�t\�z��%_(Ǟ��/��hԊJ� �	���Rʫ,�K�:<IF_b�wx7C�jְ�:��"�s2���ސ���Iw��N��ˍ���&��5�Y���^`�<j��?���`^��7d�.Ne&�OuTG(��Mj�#�Q�P!Nla�7Y�xJf�:��2eL�2�7��pЙ� ��E�X�f� ���L��Bv�TƘ]�kJ�S������&�ϴ��,�o�S��*_�-@�#e$$��/F�0!�?K4<����5�J��'�I��`	�1�0�ʄ�3&S:嵊e���.��	S�>���fR��&��C�=9�/�G�8�o��+Jonz^7�z8;���?�>�>�0�O������1�hK��>����J�D��8���|sMD�H���Z��2%	�u!�������r��3�Aԃ�tΓ��`�����L�p�CԺ!2��x�b�t ŋ��
�gk��tk���p�և3�!;��}l��������°M�Dy��y��8�Φ����L��#7�O�����F�(��Ex�F�K`���$�T��r�}y���[�VE�������`��ha���=�ZS���킄��8�1���!�)�V(�{A�5���Q�6�LN�������n�5o(��~r��O�*��|�A�K���6j�z)d�A��Ȧ��)�vP��)�-nql�P �\�/YD�hU��tj "�Yc�f�d{����	�F�
��r��-�X/��6j�N�NX$S���w�����7�P5
:+�
���%i��S"��QQ\�ā��	�v�X�G2 �ѓF5
X}Vv��,�/dY"'a-^�*�Sq�M'4j��s(�i��bM�W#T����*L7��
����[o�mVW��5���ѝ��Ip�*���!��a&�Sm����F�V^���v}�:��[����z�2W"PF�'��.�8�H��s�;Z=>(5�t�S'�2����0y��	\4��F�h8;��-�ʏ�A��G�EW)��#&�R�+�w�%<+򽹩�rla�[�e��ty��fy���H2�!vr�zh+3�N:(Ư{�a�aYD�׶�`��6��&�\>�N���t��5�9N�'9�O�CAnכ���z����ғ���l��`�i�ڶ�EZ&�c]<<���aj���`J�����F���ص*�hFh�ޫ͆�|7�ܛ�88a���A^>ԃ�Ц=��o֏�2O�Ҋ����R6>9�J���}�vkXrQ_���)��)|=yǎ��Y��r�ߤ�|�i�t	PL����"HWġ�� cV�&k��2TN��Ĳ��z��0�K��Z S�U�ï�9���\�2��i=BYLڷ��	�#����������]��Bڂ�h5���yK-�p�fظe�9����R¨������@������Hb]�j/s�����D���D-1U���q��S^�8,v���7�D��.�"/�x��� r;h�^낷��%T��r~��*�0�ͺ����""�:����ۥ�ր��u;Wy)�c_]㲍Xm`��	���uj��*�M��rX�:q�B�26i��^�ۄ�kA�FpK�(�?N��vЀ�Jk%0b��c�}�}D����Ӱ������]K$���?U�?n�>���%��tt�����<%�^�$� bˈ�Y�퉘%���;�4><�K�FឦYt9�Ϧ������x���?d�?�S�fo�O���bd��Q��>OalDK�m�l\��@K�i��hBb���Z&;
d͂w�ܡ(�ʂ�'��Qu����zs�Z�QʝD���>1�wS9�I����Byte��WLd��>�z���V�5`���7��8"M�.ڀ�1���C�.֧07ӵ��W��i&<~��.�QR�� �Bv��:��Ũ�+u=1���Bg�&��뉽��i%�x�$LP�<�7���_��
�4����X�N�:�'���j��>(��Pt1 ݝ 1R\rH��8�-��/y���I ���;�n����C`$��cB=rQ�(s�� Th�W��6J�f�wR��pV�Q>�p�<
��y�n�)�S��5B-�AQ�X�Ù�=n4c^��@XNF]h���Ĭe���v8���",[
��3�X���8��H����hV���Y$_PF+6����m���&
x04���^|~��"�bU�}�5շ�t�&�����(WX2s���>�����'h�|�*,E_>�Y�4#f�
2W9�u�Q̵ɉ{w�ݸh6����︚I�K��#��n1�e1L���"����B?���}��WjO.���ä�-&�:e��~�T@�E��1�t��M���;�'����%��i$���ͨF�|Q�t�,��/m���y�Н�I7m��d����NL.#Uh� ��#��Fgv�FNWU�����| G��i;���t BB��r�p���jE1�/�;���o:�F����R@1�7�>*��,P�9m���"%��~ q���2I����*&ڛ�?��C�}X(���XG<h1��J��������{YdB��.S�;{5��C:��
��8�(�c����Y�B@���5�Q �Q�rS��:���~�"�/?u����#�_���	˼��徒l�Z�*D�IO��6��v#�,P�gNE;�~*�o<�+̮���pe0���� nHA��M.�\��G�!G�R���6��u�Z�z->�jEJ�}1������|#� `r�����I`�cz.GA��i\�i�)"g@�G�B�f$�B��9�[@��E�T'�w{��0�R�(=�T	�:L�f���CcЈ������e�$�`rm�$Q�8�sAj0�Ȥk�1�y��y��B�}���Q�v���z�������S��T��6.�n�����X�`f&9Dkۢ��*1e���T33g�'����_��"�(  :�SDg��D��+G}�!�A�Bv�,#��_�_�`���e��=f���S/�HNU_�Q�`����"��)͏r岾y��J�h�n+���67~�Ã���Gq�����BجF�kd	�W��v=�v�*T��z<Dr������}A||��H<�lS1�ȠMt3�9�G�zJ�m�qO.�"�d���MQQ�@o�Z^���,_*���f��/˙��O�M^#}�K���ZNhq �x9�~����:T<�� ��\���	
�Ƨ�4����	1��*]Y@
������Q<!n�_�-�� ��'�_�������:"��؂�R�(��I���O���� NSa,�0���Fa�8��BgLlI�ȴ2#Y��g�U7�/�O�?W'�)� (�{ͮ�vv�f�$�I
��nC�� I.��[n����R�o��a �:oPMti���E�wp�b+�h��EL��f]-�1-����e�6�~Q�j���-�nr\�2v���o��yCmp�`�hg�&b(��κ�^�B�'i��yQ���&�^��b+�1��K�%�=���6��O��)��j��a�s�`���w��.���V1�)G������)�⁤��,]�~B7+1](�+��|%q�ՓrZIieo��n+�����ԕ�|��87_�N� �]I6��T3�ӌ�uO�m�=�ު|�B�p��s�0��o�;PWRF�/��ډ<��u�݌���Ӎ�t�s���A[��F�M��m3'>�四�8��Y�4̑�G�����q�!�aȦJ�� �U�B�*�2��u�@�82=3�ܺX��!`G̡��{XU��q�i#FnI#�T։�u{�`�"�����_ s#m�lD��"[S�6�`f�.�,���r��t�vY-����	K����S�;"+�K#����Q����H���Y�,���e�����+�?H6�d�[�?�a���C,���)Qq��a�©$��D��B��s�4;{�xE����ChM?���`U�[߄gZ��w��
;Z#Xe��J
	ܗoa|�A�f(����W����ϭN����뽝�vvQ`z�R����9>s�f�:�A�ek]��q���j��,�|��]���ߊ�.�ץ(}I6�Φ/ET����gѝ���-��ʌ�)�򂴏�L�D(�9��a�����}e{��Q��g�q)��d�Fk�1�l�����1�^��l�tF���:v` ԺȌi���y��hx�X3���A+b�a�3�m�"��b k��kM�K,w�q���אCy�p�8�$C���̼�+A���۷'��:DS�[��*���H#_3�wU� ��~b��^���x٪z����P��?w
#X�G�[�0oӏ)���9�4}���Ԍ�S,7
W| *ՠ��y�Ʋ��]����1���v7]���<Vl%n*���9+=l�9��"@�a;�e������I]����Ԙݐ��2�@wWUY͢nN.�U*�T��-%+��W�.�*���B�Xt64.�Q�Ul�63(,��,���/�{��[�a��c�MsV��3ݭ�ώ6��ſ��1�?�J~BMO�I�8����1S��@���e���ӎ�o��<�.o�t����N;]�Q�,+.	_�|�&�mU1��ċp�F��WAe�S�E�g�����E���m��p�5N�_Mu(�s���LYW�-.��9���Kݘː�>z�'�	QG�ʉ���1y���c���Ω���[n[��#!����(j�f�ISę��p��P7)Y��:\ߺ�h3�݁���^��K����C���@�Wl��!�}i�����Qmf�M_�ޤ�y�^h��9�-3����{�������:!�|dB����f#�ޜoNz�6�~��z�I���#_âNx��>4n�� �������s�^Q�!��BZ����y!�g
�:�7C�Q�%�ǵ}��j�B1��96t��n�{���d�+��-����W�p~��/�����Y�a���N�=~H�����<A^w�-#��D.0�bJT�R�G�a �j��)Ii9-wM�k��2����@�Fp~�D�F���+�;�@H��-\*I��B�o��)o+��V�N�f U��"�waѶ��ԫ���g�����q��Zx�\�Z�&	�8�I�o����%����� A�v�䢷��܎:�/����J!��ܧ��	�ɥ��1�.�h�u�3��#��"]ߝa�����k�P��尦��~��-f�Y�͂�]���/�[�n�����ݬ�x �3��.JRK�:��n���%Z�rQ ��b���f�P,�e!�w��3ܸ¹�(o.���X 
�Z";����Ʃs�Y��4��_����� ֘��1WP�d�	^OA�!�6m��p/s��3�K��ΟI�G���C����}L�f���)� }��:ҩ���NP�=��ܨ6���:�o�HNf&M��u��t��7�vO��x@CO(���x"w�2�E�k/et��\�2��0Uz������,��qd�<�+��}9���^����k�fk�,	^�[�/�Յ�5ε7�����?�syR�UުRӱ1r8v���i
4�Dҧv��)�+�is�HI�:ay7�tfF����u�}��B�+�͖�i����R�`|�R�T��/���u�{�F���-4�,�Rܦ��g����B�֗/	�c�sE��"5��PCY-�S�^�}�*��D�\�:Ĭ���D�ŇEmW���;�%��;���61cBCI�o�5���ⱬ50���$�TTS*�[9�b�N��s��nS���S+�A	O<c�:L\��K��o�8�z"l��~�'�m�e:���س���������e�>p��V�~ �ї�s^��~���|�!Wl	nЄ���3�p��R`��7/R�4hD[�2T(����;_��J$r�₞�j�91$��0T�V�nJsOr ��3�5�M�铦�ċ���/_��Y��5�P��U�#�tD�r�����BF��X���:�k���2^v��_���~�b��ƅR�0�߃�� �*��
�x)D�4��z�� :�*���F�[��F5���6�g)6c�7��jw�w�X��srWOJ�\E�R���~$�Q\����$c�b7���Qr�� ���gFe]���ܿ�;�'����u�f���P�9y㤝^�qٟ6Xl�P2uT-8��'�2x*�pV3/�7��_����DɁ��:��(H�*I=�L/�)�
�����Ҵ0~�>�VT�8�}��CVĸdL�%��ĉ��o��rg�}��8(�Ќ嘫�"w3�	�Xb��_�[�n�{�ME	>q��~���c���R���eJ�Acy��"�Q1%AI=�ȁ��-5�vp8��x]��~��˵sg�����]�d�1��rs�ե�GSZ�[��˭�ƎC�F��3�u�Ȗ����q�q˄X@���z���24��@aוF��d��|�
�����8�`"q�}3��Ȳ�M�s	 h�-���-�b�B�d����Il-Ɯ��YZ��t0~��^-���e;ԗ�٬��pW�A.���^vdYu�7^Ş��9��Y ��m>�������e�a�:�ev1��\�����=\�5�v�=y{R��k�w�)M*] �1�x��P�l \LR�N#�AWYb݋�,D
OP�qh���d�2��`I�K!O�	�m{�E���7^q�%��᭸��H����W'&P;���ua��9z��S�iI�(x��O�(^�HVa>��>���[�ibh
qlX�%^9���u.�#m�f	d�0ƞ��\�P&/5z9��l�0d��1�5�I�ȵ�5���� 9� ��ͪe&�7b��C��|�g7f�5��c���Bq�T[F{�:I�s��D� �s�L48��r��o>�O~#%=w��fk�esH�?{�9Q�UFn�/	E �<�lW����O�6�K�u���a��3"��vl����=5(ӛZ߹S�����~�%l�ʪ]�C��@ <���f�t�����p�����+�K���K�J����3���$�D���y�A��M��P�z�KT\;0�rDTo�d��m��=s���@�}�_;qQk�SKD�_wR�+� =�:�lI؀���T1�G�����&����������T��$.u���i��&�zv���
�fv��D�vB�i�}d�?�I���'������t&���!'��%�Ϋs��Wg�[i:�����;��^;��74��&
Mс}!�-���\�7��vW��Պ��,n�*X�:�K(�u�俨k�;mG�s�LC	�CNNe����g�Gf1�\I�Wx+Sc���9�#�F��`͔� I�� �4J���VZ"rv�������������
<���ͳ�z���[�H�A��{}���އ�Q�$F�V�'��"G����9�=&0�z:�3wɭ[�sݽk	1�B��z;�FaR�n�D�{��r2�jo-��+3�>��#i%���1@���ѳ���5<^��scJ���G��f�&&09�R��������nC8�T�1%@���S�bI�3f4H����{�,�=����+[i[L��k;��ա����&SŢ������N�#vH}Ʋ�x=,��=���$���mMl���M�KR�ӎ�u��UV�t�h�X�07�(�K���K��V�����;:����؆W�aV�=Y\5`��]:�g��3�0g�+u��g�M��K� ��U\��\WkШu���/#�Q�aa�Y���)0��K�%�^%�X���W:>�چ�5e6n�M���'�+8O��N�C��p��z��e.:vaR2�c�=����Ѝ���]��X<�vr赓�&-
 I�X`NI�jS���)7��q����<�Zr��0_���	B��"�Ҹx�(�`���}���&�0�'W��h�6G���1/-��DB��]zyn�w�����2}��O����][�������h"���N@9���� n 8ݩ"I�>�Ld�6H�׆��7t�p�D��š1�"0��c7m��ϖ��Z uY���P^���0�?+ X[�����u�ߢ�a\X�]�{g]��vj�O�	���[�f%��s!�
�|ʯs,/}�ۻ��2��MFO�,��.O�s~a;�-��ڃ^�X���\�qغJ��(�^=�QyL�ݎ�k������bd�i���X���D�� #�"������ ��F]��x�\Û{�t�1�ǥ�諭�Y�f:�ƹ��m�F��[	p�#�Le;��Ą6�46!Y�0uu-�|$4���=�n�=�ȌY#���1�Wy��t8 ��t7�#�ad�H���(�������K���5M��C�i��4�荀��]�o�jJ�n�
�j942�t��`�-օCJ
"+������/Ӥ�ϒ�BE��E�Bʤ�0:�%:A>�m��Q�C��@�?�@jü�Egn�� ۲ַ{<�rgϨ$�M���6Y�/UР����;����FV1��QBJNO}dO+ۘ�m[Ί�S���a�U<f�|
��1�*�+."��G�dp�+P$7�u�>Y�i���D�\�}w^z
��
o���5DY�1!������|
��fC���i��v
N���:^�U�9�cO8�C�o��9����ƫ��䓍a޶H�EumǊ��YQ���@7\����Xr�bm�a�vca�P�*DKV"qvt�s'� O%�c=S$�Q�,�;�k�{�"���ˁ�ܿr/gt2�xJn4AԺcȁT�tR�CξC�b��b�.Qf5QU���D%�v˽���?��0�Eb�aJs?�N2�hq����i�{c1�MEU����)�|��{%��0�9������
a�*�����!:C]��3zC�'V�L��k]��
�{+��G� j�I�}#��l;��o��?^I�RGZI�D���z��l;��$���x�rX��Ӌ!#w�[�$�=i���JWh�N%6PG��M��w�'g�����-��AQ���4��6����-��Җ�	o�49eW���-2Y��!�}=�����`}�	�����{_���rU�S�Sv�4��H{�HR���ke��c���E(�n�_�f<u�>�	�تX������`P��oVk8v�����jkP6*��j;�ʿ�&~d���_oIH�m���%>RY����.sT�!�I���2�� � S��
��yM�g"o����4���@�y)���uR�LeL[0���/ T'd��XT�*�����e�����&s��✫�J�"8����Ѩ����ǆg��T��DT���h�ةK8�� �VH���KI��շ,e���RWK�U���A�`�Ml�����jO�5�ɢxByBhͧ |�������aH0?N���᪨'h3�`�@��<�����ND8���G��$�v�&�O�W-w��?8��з�`��9�����˝�D�6�.xcڣ�=��/��t'��6�&h�*(��֚�e��f�"��AF`��%�,o������#���y��
m�[
��L3_�KF��QOZ[�����K![b�_w�onq2�#\�tm��g��C����q�V�*"��X�iQu�����T嬪�K�v��r���n/@����7� R�X%��D|�_� WPH���gִ�q�i�a
�0���c%b���ܟ3_eٴJ��O� ����Q���i� �ڜr�[����{Uq&�����-��7���p��T��э/8�-}�x�!���V`�r6� ��{��S��f.tt��ƈ���W������W�Ʀ�lg�-�q�'��?tMi��
���Ph�ݖ�7���L����|�$~.�9���b0p�Xp�j���^Ơ�\ȯ��(A�"��v���,]<:�C��B�P���b;x�#+zv���4x>F�K�=�@1n���TZ4�����ɏ��J>8�����G�8Wũ�<D</3��r�ENV��-Y_��}�i�+�2\���}���l���l������4ؘ��%�3�\��s�(��4��Q����6z�X]2@l�G�p�"GqD�@��_ʜ�%��r6RA(�轼}��k��WL��C�`F�5
�����}���ZL&���)&�8�*�$�Gֽ^�������F92>�4HɅr�nnZw4��AЉ���ʩ|������m���J咒�v��Z�2�M�{ӛt�����5�C=�I%��Б�lv�ml��3�͝���]�L��{&�hw�����P�f�O�NL�׊��)��\��� B
W���)[����/9�����+BΘ8�7�Q;A�!�%���ä����n���}���]�r@~�^f��3(�u���>�g3-�3B2�"'I�����\Qq{p#�p�K	�7�TŴ�۩o�=�������Z�y5�Ty��W�8����4����<��"S�!xX��H'`EA�U���]��:W-�R�1"��>^4����g1yo��4mi����6������u�����fL�]�|)���I���-I�\TVO���z[{��X�u�ʻK�>�p�x����WU'�]#Z�� ĕm(C��K0�d$�^7ELj.��j��_���7K`�H�40� d�x4�x4���ϲ�
����j�v���|�=ڌ4Q/�#+Y��s���]R�Z���vA��b�a8�ΪRb�^,�.�����/�a�G�5���Z�k�,�y�!RP�����N�0����)�Kx0�Ɔ
��H%J�]�YW�7`!�/�6C�#bu#�y++{���Lps0���Э|X���ݾS�{����X!�ݏJK[�TJ���xi^2~#/V��#��]����kwg�_�.�����&�*��Y/�_��h
�D�	cE9�%��6~%�����DF��]��#X0�K��_�7�{;f+���	-�qe�q��mb�w�B]Ӱ=�=\�����&���6h��?5X`8t ����=Q�]��(�u�v��V��wt�����S�����|��P߽���CfbP�7:��x�{܇��K1�:G��:�q:�21�N���|�4x'��q�բ��d�X�<C����Cy@b\��в�J���wG+q��r^���fLHև��;H}��d����LU�9J�YN[K)�X�#�g�]']ws��td}�*�Ud�{�п�����N���%�#Fm'���);s՝�p�A,�üX"��r�Ź*m�f=��	��;��$b[�����|W4��l��I�0Cmg�g��J��n���hX]�ӻ��)[�-��>+A���������@�5Q|��4|�V+�v��{[6�0��K�r�^��?�n%{{?{(� 32�	-�AyQ���d"1}��l�7�Ӝ�?�v�9]r:�U*��_��T������OFVݴ+���l`m���ڇP��A
��M� @���p���%�z�Ћ@�8;���7�@Gݬ�@ZkӋ�������1��(����E[w��/�ԃց�{r:��8�.ߠ�$�<x-~�u�9��Q�R�C�-���$p:=_RԌ�����h���a�вw�N�Old�|���(5b�	�B�,��p�A�H	]Mo;��w�>q�����X%����=�S ���`	��ʟjK�9�K5������^���������I?�^��"&���:�(��^=+i��H��cͷ��P�a�_�m�:=�o�8ވ����H)�"��>��Y�����aw���:"��o[㦜���	�bw4r&�i��ݒ���Зbq�����ٿӢ5�8�1����ʨxW�%�L�k@(4��OlkIo�	i�	���W1���p-b�g,iw�Y�Ae�'��SC����ƅla�MX�-|��2O�W�C9Tͱ{�{�_��H�c���S+(�%��r[��&��<��/����f5ɬ�#�����<�.�E�=\��9��9����jL}M_ܧ
lg��E�N�7S�v=�]��cL���^��2q��p�����g{�PC�	�1ܖ�A����f�;~���gBSշ��qW����JQ:�(B��a�;1�6C;�� S����5��j��`} �B���9-v�#�.w�Y\���ӿ�h
��s���� 
�x�h��07���W�T2y~�m>��P�.ܭ���*	��|-,�l�PgNq�D8����\7�7��z��_�S(���]{�6�vS�M���.P���ʽ��ǵ]9C�/���W7㒂�Cdu
�9�n�Ȅ{����s��F6Ǚ)�,D��U��7%�hH�(ԏ	؞������M�����W��j蛼y�Ĵu�i�H'�´v��P�gxsӮхȹ����5z���P��~��u�6�W���?��Jtڀu�T�(����2��F�'�5=l.(Wӌ�N?���Fp�������D�� �^�)9����F*������i�����m�������z��x���丟p�Y Q�q��%%�@���^��)�0� ��Ly9Y�9&Aq�3�����` �v�e�����a���	��ԫq�l����������m��Z@ȏ2l�ƗӨX��c�lo��q~���~���C���uF���je�G��d���~������xF���.o�,����hò#�����$/�KT��i���f��R����D��Y=�"G,E�op`���"�0i��_/�|w���	��{�r�Y���W����W\MQꖽ���g�԰&}�ɉ�4���i%���trQ�0���	0H����(6'c�F��,�g��8(>ZR�qڽ7��k$^V��#��a�8\a��r����1��}��ߤ/�߸<⁁P#�Z��w�yW���
��c�QmwR�PJ?jlRC�}��	M��@bK�`��µ�Y-Pܨ�15��wwE8C8��Q:&޻͙��o��n'��h�Ѩ�AV ��4����1j�vǙ��3q���|
$`b���B����8� �.��'j㕦.��.e;�|��8�|5A����KA�qxD��*:����he�ժ�'*C�(n���"���c���Xt�SS�f�Re$#kˮ=�++�p��B���!�9!?X�.�&m��Q�R) T���nf�'�M��׾ӭ%ҟ�1#ٸ�D�#mأ݇H��'�o'\�bd��1�6�Y��_ ?A
���D��b��1���܄�,�|��3��B!/�����(�����M���?������<uᅸm.��̟�|�^�O*�z5�2�E��:�>Y0�q2�,"��*iR0��s���6MS�� ��&:��M@k�uē�|�Q����?���Wg�ق����ې5���j5���넙�Fbx" Vg̒!C�� ���d_�"�r�m:�B�=?N�&���=�9Wך6�=� ���{g��{5����V0�w�������|�/�2�Ϡ��;V�ק�Ft֖�c9k��f\(�~�,T;`�� 1pV@�E��9�9�,����t<�f�0�ߜi~xt��� ��\���+g=g��c�S�\ܟl(�__Y>��Y�I�`���r���+�y6r\� WsVT�t������q�!멂�H��Y���pmK�eP-^D�8�s�}���~N߽�5��Ê�PQ������)ވ��"w�d�ioc���g=ox�N%J�.A0#5��n��U�i��f�MT�<(�(_Wכ-�����)|�f��E��[���(�����+�>�)j2��y�tM/���d��R|�$���M��'Zj��,�^i�/��C�˄�<�foZQ����U�n���?r��ū�'Ǖ-��!�vd��t�
���R� ��	��|(t��BH >�55`� ��8�؊�$:2�2]�3?d��#�o����d���v�ФB�h��]��5Qb)�Q{F�ބ�pԘ�IS�d]ıu"��}�a nK�	!�g�o��}�N� �؞E�
�0�;�T�y*A��X \;�읚��N��e�)f�S�{�.��u��ݻT������T��Xn���P&�N�C�����=̄C7b$>p�L�FG���5q����������%#�g��ƀ�w~���m�j���U�Bu��.�V��G@��ɏ��ah1E�z�В�h,~�m����+	������]�{NXe[��; �Ceg�3y(�I1L��
� �h��7Q-��/2���׸Ȥ�>g�4�a��,���I�%�����):�E&��O�GJ��e|a����fZ��m���⪜#����1d�8��=�����m㡹!����f�g��~n9X�	TȹU(곱�(�,�^��1ߣ��	)!��(7�Y��ڜn:JKS+�@��"�4�ǰ�@�6��1g5��%v
^��Ԏ�*��Phh�\�����?�W�
�1�R�� |�u��
_KKyy�j��{�8-졵D!�r��rb�8�#��Ξ�l���{�6�2�c����_�N�q0�G�oChh����m���Li�؍S6|����E�c�����ώ��cB�7�L���B	E�XHR�X_��ޥ�#�mibf�d�e�1���)�^ &O�Fܮ������ӵ����z���R2H/2�SDm'3夕|�����s�O��9�xv��0r�X���;��L+�?���qfk�A0��׳�D0c1,��4�~�h@�f��p2��)Ԣj%���x��Jlל1%d9�)����q���)E��M���t��[Z����w�|^2��pk������ZI�l+N"��mw��G�EĖw���?�c=#ha����JV�;��F:d�ђ�m|/9%��v��zY�s)ɉ3i�f^�)�>�'h6�C'��I��o�:��G3:�b=A���"��a��s�B]��0[C/�/Ҋ���ł��	�������?����.�02!C��#��]��ƙI>�n0NBp��V�[�Z�n2����VN鏘	�>xJ��Lp�%3_PE2��j��UF\R�� �4N�g<�5�����,9$0��a�c��ܙŲ{��\5}��ƴ���"�|G���	�Q��1U�3�3�|��,J9L�ڽ��������ZR�l�W��"�jY���1�]<0�J"�E�/����gU���D�D#�����Æ �p&��0>��IT����t���ouj��B�\�����no=�C)���/4n�	��0�P/��ŵs"�5�W�W�S�9yC*�xE��C�uG�JX�d^m��b�� d:l�B�xE������DX&�W����1�]w(�P|��!��Ġ�ћ��	|6���<L>������A�q�C+�2��g{YF�n)o+f��I��/~�R ��8L���^3�#׊ю�ç���I�=D��r8��(�S���«���ե���_����_MO<ySR U���P��8��H!�:�y2��$e������O��N?
��*�"�]��w\�ˌ(�az#e����ܴ-|5�Sy�\���U����l}*��e3��p������	 fJHj��L`Ϫ�[ի��2\T��RFi��X	zY����Π�t�C��Ș"z�݈NV�`�j����AX� 2q���+��X���a#8N�c�Xc"�|�4\��_7�!	Ų�W ���=�Nk��`�D43���QF�3^��r`?f��Dw=D�7QPNO_U,�
f�ĵ���i=�'�X�ɀ��9�����Jf�թ�f'�t�_|܃��d|69Ͽ��z�C������
t[���T��3S�=:&�
�֒K�BOC�ro�,Z�4����Y�{�~g�M�FL�q�3�m�9w���;:{
m��.�m/��X���R�.�����W�����^u�������<�b�l�9���R��j<��_�+U
�(�¿����{��t@oom^��M�J�H�>����e�Z �.��ʯ�,%�e�Yq��"_������9wx<fg�
�����xٚ�E9,�$�0C�g3 ��c�&���?v�F�$Q	�����;���R�[J�/�I��ӓ@��4�(-�I��o���<g�%N�6��>� ޕ�p����Rc�8V�	l�<�a/���kK�j�)��Z��g��}p����0�]ޣ�Y��Lps0>�8�^�!��lBä�P}����?����)}�������Q�- ��v��r��b�ݍΐ+�F��p i���m����+aZVc$B�J�Y�mr�rأ���[�?l.��VZ�&���<)6" ��� �Ze'�n+�G���_/ަD6�������37��/��A�׸�Ky�}$�D���ޭC.f�z��\�2H�xC��hP�Ni�ys4L�T�`�OQ*��)��`O�)`B�9�7.,���Q��hf��/ǹ�)|�K&�t1��@����	~��a��ݨy����b��s�m!�
Ѓ�1����l��1aCq]a��A4���l�.���T4�t����S�;Ԝ���謹�_��6�p�?�԰t��� T�b��l!��V���)�c�#�����J�lҿ�O-������<W����u�&3S�h������ѷ�o5�
�4�Y�.h��ǕL�8$^ �k0�}�i�1!�Bb�pt� ����%r_���P�$&�D����m4���/�n%��k��P�'g
5�H�Ǐ�q(r��-ϕ���7L�#z��(Rk~@�|:�:��#B@���9SZm�Gu�E�ȷ�U�nB��j����0Ç���*&�����A�"A�1�n*��})��,�irC	l��y��g{n�owm��Kq���}����ۈ�ua��.xዛ�w�r�����w	W���i���)?�w�F�Zؿ��Xj��*��������)���2�P?��ඟ�o���q�Lv����Q�#�Z^�>9�}>ѭC�\m ��O�׬�W߾-Q���kn׈)�ڣ#⎠�z�7��w/�9^r	�폯�nH��2���;֏�Α�LcHֻ�	'���S�}��9T�k"���`����)m��	�kqX���c�6+ey��A&��<�lh�p�T+[*��c��������!�����4�1ќ��*ڒؤ���s��mO�1}�HcXLʮ7Фº^�B�Խ�����<yR�ob �ê���l7����i���h�:��F�7�`6��%��4+}�Y7�A&�Ed5O���'�"q��R��Z������9Rmخ�jw1�������Qw��\���:}u�H+�����aGD$	�Xe��`�e찏#C�G���B�GЩ]���IUf��@��$���"(��.[�7�ϯm�F��	�ٱ���}܀�g��ͺM�~���2��)oȰ[+���y���lf~J��|���=ˍ3�A06�>R>7����ۈ�bY�Tc%k�^d�j)�ꂊ�&p�����
J�=�d�v�d۽)"9f�@�l`�*%�d��#��ԍ���s%RՄ�^T�~��O�ṃ�N���l���1D*���aq�v�a����01� �l�Wԥa���0�U�f{��83.��5�f�"��ѫ�ʥ��(�U+�Ǐ���+�1	7�c��W���T̅�qȉ�:�j�C��q0cjW�#?��[��Y�ӿ	x���f7�l1�-�,m4L5��-RN(������eI����gs��&�שƢ'go�_�v��`M�h*�b(�$]����.�8�X����J?y��~��4�ZΏ��=>>����&ޖ��^*��K��G�%���;��1 ����cɪ�3i!���z��^G.+�r��]W�y�� �wC����7ƺ�"�|�ȹ?�l�\�(�����X��S�C��p����ǅ͠��.�V��[K���ކ��
!��� g03��'f����I�I�j�b��-�U�`�7����@��=�~�U�k^�p��I?%����᫇�O�|��$�x��c�y"`FW z`s�htsD�GUd�D��`툐)3����{t+xQ��TB�w�`��S�6��G��^f�>��[��E����y��Mt������;�BXn�F��Ѷ� �n���J��_�#ъ'�e""�iA���|���n' ��%t/�ms��׶��
A-��]p�<�/ɭ}0[$-&�6!;��{�A~���+T�09B�!:U-�f�r4��
�"�K=\����i�H���@��f<�vs":0�Dd-��f�Vt_2�g�u��G�w½^����v����g=���Z��s:�߃�1���ԍAx���������c$5ô<��y��մ�@;�C5^�_�r�mu�$d��:%76���	EqǮ�J�;=������ph���'l����Z��:��24҃��b�o��)��-992�5	�̬�����w�Z&4��i�h���E��F����+i��q'�g��}�Y݁E6���-�YǬoX�zj;�|) �'�Ҙ��z�c�E��=��z.��2�1�՚�:���k�4<�;Q��U�H;u���v�'N��&ʠ���|��(
�
y�$���Wc^ټ�<�Xn|p�>af+;�μ�K��&�d��{-O-7wKٮGFW7�����a�H�Ux���bn��j6.B��*��V��nf;:�280 �C���w!����O���#���⃨����K*�&�d��J0��Y˫(�R��ч�Y�t=�b��{��K����.�.�:c%O]9Gp�2�Q�69���EZ%T(e�M�7��J:e�C9�@*�敮�����j`�3? +$ 8�0�|�i��O��ƒ}"��4o���H�B0���8��X�O�5Dg��}Un���[QWGJ�|N��¦�������-��T����S��e�Rp��%�0��]�Cfu����5ȐtرcWvsIJrT���I���4�9gV�܅5�oWg�r�47���a��ݔuMQc��l�8�YC3Of��C�4�wf9�y��g�)%���ލ6�Q� 	�G�DWJ��+iRl@��%S������KT�#�}|��,��ת���Q;���0��
��.�6��5�̄�e����/B�nR��;���f�F���p��m�w3���#�X��F�!U����(I`�h�}9W�Ol<w�E�
Gl'`:���(�"y�ՙR!T)�T"�9i=�@ya�<�� 5�L��]�p9cR�u�&�!O���V�V6���`s�$���N�,.Z��ԋ�a��)JV�.�Z_熻���֏�#s��<���5�B��Jjt�Hu�,Q������`��<���>�?'P|�T(�D4��:�0����?;84��p#ϡi���4����Ck�)J��/sW=I��Ww�aߓ��_3���	����h��^���V*�j`2�Hp�@?�
�&�������FX����]fh���9Sb!i=u)'���N�Wh�����ǜ���\��?���N�T�!��. �ؒ��_h���@q��8�$y��|$d���ԮF�nUHE=��D�@K+Fo�zI��L�p	�ID �&�L����,juۺO�u���X�l�Zc�:B��Ò�5_��{G��Z���VĄi�(�i�F��M�DA�z�^җG��1z�aQ8.��5c���k�}mG)
���<�+�e���'�de	�sU�Tv���6�֤صh:��~]� m�8Is�dDZo ���DL+t��m�J�~x��U��%��)��W������ ���9h!ƹ'��#��=�x�,�P����y+/��Ynm6HԳ:G�{s���%d_��u<�C�D1O��㎹!π�v5Pͩao�S�]��!O�A�< >;��\��_՘��eR����hh�b�W4���Wtj5�P8�O_�i+��#F8Km�QϼzM� c-*�T�6������ɿe)P/|}4�֢Cݒ&g�Cg�$U�	c�ҵ��,r�!�@�;z����v��[<h��k�h�MnҜ经U���\y�W�J�ÿr�Tg�?'��z�βpkdic�]
 Y�!�O��~��H�`DOw?�HhW@:uԔj�%�Բ�M�`�}���	�uol[����/��o蓥9���V��bu�a.��H�Xc�d�j6ي�dUċ��5���_%�A��[��[/��D�SW�~77ꅱ�p��P8z���ޛ|�*����'�(8sYSB�.���Ic܄{�`_��ZE����?4��a�^v:
�oH�L�;k�v�g,�P������k��E�w�'�D��9��ĩ��r9��O��=�X,������E<�:5�n�|�
��P��K)�A%�=S�13��TP���r].j����g�$�Un��~Z&���V[F���_N�E����D�ķ3�^ca4�T��E�C����I����U='��s�#Y���v��ލ�onÞ��xxV�ܣ�XW|���頚q�^�\2R����d�ː�t:Zf/���Mƥ��UC�+�t^q<^�pYg���:��Bn�}%i�IN*B�CA�J�I%iǁ�l���f�Xf�/H�$�1M��/���f�Q cn�U��Ӄpe�(����'?Q$��N�6������獫��A���/	p���w�6����d��

$�Xr��[���W7��`30Δ��.46N�&֥�V�}�f���q�k�幣Y�#�f�?��mȶ���A��$�| ?Q�G?vʞ�j�P��3��Ʌ ����-&��?a��H�����\���#~)D��0��.%4������/~:ǱO�9p�,7�÷d�iX���w&�-Utգ�s��_����2�h��؋@�RC�Ŷ)87��Ű�H�l��:��@�[jU\��i�g�J.�x�l�&��$���Ax׻��Xsd���>���{`!o��Fqq���q�#�s�5(/�ْA����2�s�����r9AB�n&�#������\"�&��ʡ1�o�|�8��4�M5����؉!i�#
�ё�(�x�B�h��O�����2 W�U�3J��/�|)B��?7�n�[D˨����!/�?5�V9���CY{��$Y��'�p����-�z	��D��R	�k��-t5x�J��\�E���p��Lka:(�c�7����� �E맴¨���tm�bj[ة�IM���];u�A��k�p����=Tg�=��%�=��P�)�Χ��6��$�"��K��4]>vXߔ�����>�Y'Bb(+�s袏��eo-b�e^R���M�N��u�LS������*����nm�G���KS4w^��Q� ��8�qY=Y\7�	����X�{��+;�ӝ�����^J�8=d�f	�`LN��R��#7v���J���f}����U�ؖKY`e�{^�4�םơ�m\Nc�49� /�w�X��u��Ⱦ��[<[2>�n�����[(ʟ��F����[���O����^V��+݈:���Knf�TC]r,�Kͨ�=b3�)����PenQy��n��UOt���-Y1l�!�*��}ݒ���v13u�dw�� �|�Ru��F�A��v�P�p�@�����E]�
���mw��?��,�-V}�PG-��*�?�?��Ç'�,�b��c�����%y��>t���C�P%���*�|#��,���f�k���j���)�� ?I�=���&ɡ��{<�юKCW򶀷�a}��݅=��{�kK���Ch��C�Y�M��Ŧ�0�=�����d������,�F�v���0�a=E�Fĺp܊!�=�_��I�iI��V��nR�=��s��ӓ�e�C����mV$��I�T�\W����nw!�Ws�	��En���5����jB�*�|��*v�j���e���x��$���ȶ��0���")��G���Y���:�M닇O(��I�ޔ^<* �7$�@r�di�;%�gs��r��X4�wV���2p�8�>��!�'�K�����GW�_���`AO3����p>;~PV�D�馊�t��Cаc��gx�t�Vu����r�p�VQfݫABC�;�	*�mI�>�P����.&�������J��י�8�izEa��`�.}޷�W)Ӳ�� ��cdq�>�־���zY����y�E�3'8��8�N籄E	�A��C<vc\5���	��<�߈��I%��t��J��A���V�,Ŕ�:"�t��b��e����(<���2��o1�O��	7��:�ՑD7�*yF"յ�[�;�)��eJ�G����[ԛ�a���V��[�>�0;��5e�'^��Y+'��#5i9���հ����.r��*[�{�x��7m���W������H�lLʋQ��N$�1E�M*O�2]�H��uA�ƫ
8`��yRB���Yj~ۗ.��<�n��6�}�gjO&fz#�~�F���ނo���� ���>��s���l\t��A�b�c���B پX_�B���T'�S�s1Nx���X1B,�_��{��7���'^�kp��ӷ���5�M���&%�i�Շ��;��1X(��J���v��c�FN1Ʀ��� ���%�̸����A�Qh����D�{��t��2R����I�I�rd�ˇ�q2O;�V���%�'�FlF��{֔KJ"�� �ݙ9Ċ�#�f��y��{��;�6�DR\�C��U6~��--��s1=V{4p�A��5�*���Hf�pN�P�"�hQ�t|��]m?A��߁�Z��Gyּ��C�SlEDQ�R�,�������B�.�V����w��x�+5�6��z���ڋ�|���y�%���ۂ[�%�����t��.r5�S�Q�-�N&��!��tq����'���Q��a��\�(0}�@�n�Q�I֌��g�����:s�n�Y?J���3�1�[�$ک	/��nn�� �Ulc{��� _��V��SK��_����s�pd:��^w4����䏟n�p�]T،.T�E�rN�f��P{)�p��D�]��&��Zܪ��WtʋN{�0H��?�-y1$-���k쀽X�c/'��4ƹ������\���=��ѡq������5�r�O��A;VM��s�gw�k�dsiP�Z)wl�$�\\��Y����x�M�,��땫���9t/Ņ�e�P���8.��W'H��\����bf�#�_r�nc=݄���}��Q�r���SN�F��
�%��E@�v6���<�U�C����} �ܜi�d�D&V?HZ}�G]��ꁬ���M�?��3��+�-�b5�;#��ŌT�fU�6��c�FS�yo�Z�^1CW�n��u�HG�r�X"�)Z�jL�;���Sb�F�q���Z�ٽ�T�f���s�^��oo��:�Y�B؈���#��$��~Z�	������/J���<��~'��=l$�O��"�uHg r�"޸�:<r���z�Y,�D�h~@�Z
6ճH��S4=��gmE�l=v�	��̭ r�K���L �	u�\��fC
s9b$��;���[�
|��(�0{}��2F��c>y��!�8>"��ٕ��f����}��H�#�* ' ����Ů�d��
RPҽd>X��j�;�ZV�;�;%�6�t��������4��%��e���(EJc�$�ͼR�@ÿ�G`�Uh隆���ܳ�g
�T���?����`���q�	���)m�����G�\�&���V-��0ńڂ� �M�t�6L<�)@4�.������s��M�Uˁ9��79��Oks�VukT|;�;�B�m��W�њp#�u�h���\�]�@2��S屡���,z�_��� �vVD�@ X��#��nJ6�!��[J�shڋ�p�X4�����R\)A��]m�.��m�(J)��d�ʷ��AV!��	B�b�ʥğ�L7�SI�Du!E���Ĭ����@��im��)qo���0���x5N �*���T7^� ����ez�h���s�,T�*F�B9#����@�y-d]	/���݃��k ;�q�
����1��l�b��|9���.Y$�p�/DV�ՕH��[]â,����Y{-��L���$������%���]'u��O�����%��)@� �ؖc�]��c���d_#i�\��w��kn�����v!�D�ZGe��Td���u�%1<����>�������㓉9��y~~H'wt�|Fhd����X'��76rϦ�{��v��^G!�����H϶,�r�8屴��m�9�ڐkNL��QЈj�(T�Dy.�
$�q�<^������2�ҽ�މ+A���)�❈��CA��@@�(Q���	�Į����[mʫ�������_��aqwQ�;qOvޜ�����Ì��8a�ht� �4wzU��\y����!�� �P�6yC��Ḙ��d��"�mә�������0nU���u�rà�剭*O	?���K-3L�Lv[��{�!��2p�+�돂���"	-n���!��EBO=�!Y k1�Y�	�-��X�3o�D��{�Md�*4�K!����V�6�=��1��L%QBef�;�Rs���	- ��rE9M�Z�e #�ځ�������L�ܢo���@��>W��n�0�n�z��/��Rڰ��1Q���O�٩��a�����M��[�x�#���D���6.�{,r���i~�1��\v��g܋���5�������7�~iǕ�R<�����D���-o���h;�$x�f�lQF	�eN������ CB�y&��6�[k���Jn�6��< &o��%�S�J_y��p�煅vl�����Z)	��[?����?/ީ��մԏ�Ɉ��ix�����bZ�XE���r������+_�*��2�}`�y����&��dsV�X��:V�!�K�\8{Üz�T���h#���t�眦)?�+i<�+j��A��}t|Pg�Y@�I�+9D)$�={�f2W�LEg9�Rޠ%��m�{��F7�7R41k۔hd��"���Z�.{:�w�g�dT-S�E��z5~3OCON{�Aвr�;)3D�\�����:1Jz�ly�Y]�$T��M_�3�.Q6�tK��7&�lA.%�&�LH��+nk�g��� �ʆg��0��W������ނ*K���!���R�S�/<?�P�\�=N4[�
��NM'�!�,�XW9́;�#,���Vd���b�Z��k�\�T�T+t|oCL��H|ۣ��S0�s��"���"\�~(�4]�KZR�%(e�.������H&�V���w�`ȣ�9��Y%X	���v�Y���-'xT�E4j-L-���N.����-���y�^2���*�/�DS|G�|�k�uj�	Zn���z�PtM�ŋ+�nC��6�:�.l!PK��,M��m���1�*�
�f%���Z^r>�Lygyld�[v8~!&#�k��G�k�]z�~�݄4b:�1�Y񭘫���x�N�������roև�`��[��0L�ϧ+�Ǫ�b*�a��ў�Z��q�v���i&#�Z��D��t,�v���ɔw�E0x�:#{�҇2�p�n¨���2E�$7�e՞�����&���S�"�oT��4&��$"�'ҋ�E�I���Ƞ�r�������bB���w)�{��*���J�#wײ��U��O^(<Y4u�D�b,�3�-����+�{J@ʲBTf���Y�E��A�u�0��9���!�{b�+8\�;ܸ����ߞ������@;Q���e7�����PqN�t���ڵ�DǊ��A6�G5w�W+Z�s�����/Y7LRۢ.r���j-�.�J��k��!��<�v���/'Cv����"¸S�cY���Vo�]����|�)D���;{�m5�o�?�|�A��j��f����U$=nT���eg0e�9�����p)n��a8B޿]u��=�0f<r���m�.�c5rɚiE�������2��|5{��is-� ��DK��>���1�{�K��=�˺��ů�Qӌ���TV"\���6��ܾ��u���9.��e)�;�X�m�c�jnP#.oo�@����%m���	/�)�^ϙ6?�� �B
F|�ql��L!~|L������!�c����w M�N�Ҝ�׻��\("�˨*b�!���c��E>C����Y��z��#�K��Yc������Dl!%���0~񃾹
x�v$�7�Η�Mڳ��D��b�%~=��48۬J�	=�wޯ�=�.8U�}$~h���+�מs��8��!����L�8�~���O!YE1�����bJ�O�`����\�����^~�Gcb����zEC\BK���ޖA
��UVG�%]���
;��%_�ea���d�!+��ӝ �dD:�c{Ƣ5�Ƙ��m,,��C㍧�DSYa���'(�6Q-1�Fj���JL,��y0�D3j���MQ�H��+�d����d��
���j���F��|S��nQ�h%H!�"�?2SaٟAּÔ�/����\�ZV����H�$E^�m�h�+��\��/dV���n鈚�I�G`���C:�ܕ����h��z��{ׇٺ �c�y2��@B���y��X��l>Ε�X����,W��F��<K\f�M�b�RG/9{P+#�����#�% �/N��@Co��<PTBGRoW9�q� �E����DW~8����n*��#D�]�r'~�0}���E��8�6`k�tN���!PXR�_����JN����rv�	�7�5&�-�R�H��1�~�����Icp�%৸U~��!�'�]�:(?(e{� ��m��'C%@��4E�լTPcm�Ft���X�ʣ��u�9�1�x��A�~�kE�5H|�S��Le5�܋�d��W:?T��^��2������̉��˙�֢:}?	Y��?�I�x���k[t��-�@{R��>G����J�g����ɕI�U9(���B�S�]��I+��rr=�%�p�0f.�8v��\�^���8���p����
8��FY��.����[=��������_|lM�2������@�-��98�AZ�6(2#L�+%zi��gtH��Y��~v��Y)�sʠةs|�F��MS-�����h&���W`�nŧ�ۥe\�C�c���G��`�ZM6zIlYtXe�h,�� ��[�;6�!�U��>Н����������'�K�rH
b�a�f�9��.�G��)�"��x\����Z���\���:�2_�J�97Q�����/ �-�&�8�P���V6Agw�H;:B�u�ZQv1���~�I[�o\t�ڦOY��ʤ�lw6����P�~�h.N;m{���)��<���S(!i���M���I�b nFP��Hd�N����E���	�H3s7ir���\\ƃ D��<��0+)��h�I]�688^�j{A����+��N�(�|�!6� ͔y^��P�R��������]�'ޤ�2�[���@�-1|JLJ�)�o3�_���suP��ͤ�>q�<K����D~��#]�6�S�ĊK�����|��
u���c��La���|���0��$9x�q��'D3��R[3�!�;�mM����y��K��Y> ��R���4U���Q�[
���*�1⏬������MuD��5d=.���B�xyo���}�rMu��q�x�*�ߗ���ٙ��|+Q��F�r+���89땐��BR$&+dC>r�4�J��&�����Vf��?�!�*�b0���Id�5X� �O�՚�&�#(-�ߥ��p�Q�B%r�5}��:�3\Fj�[�C�]?�Uy�p��g�K���!��/�k�%ޱϴW�m�\R0O?'�ȇWsZ>� 8���SM��w� Kڢ
���oF�Ff	w�9&�6g[�xg�pGK�"yb�yv����vaȁ]�!o�|^��ie��!o�׳j~�as3�T�`LL8Bsv�<p�T�TC�OL�"�G��|�"�K=�2lCRhG�S��M�ŏ��),�{��(3DI�3bT>:I�{���5�
��o֐��n?�K>��"��P���@b�P�_s��Sp�G�n+8�3��:����{�dR��Q	��k4�d��D��9�C�|UT�og�U7���9}v4k�A�Ph�$���t�$m�?l��������SX�����)�k�h�Jk�����Ix��I�"�GЎ��6j �>N�Ϊ��,���U;@[��i�o
0�[POf����L��� $衃i�$=+"4�)A���Y>�Q���\���'9qq.,q�ڈ�T�1����|=ڎ�����!z|M4��`�D��C%^x��vA�`Q1xr�q6�e	x7�b��D�]�=�v�Ά��+��`L�3LɆ����w>���^��d�UR��Jt �!���� �' q6��Xy%��:.��0t�,��W�lZ��z<�Kt��;?~}��$>��n�d�l���r��/θA��UW�;Ӳ��]J�#�7Ub�����h��J1,mHGTñ��WCc�4����/�#y����Iߧ�7D��	���W���\�M{S,���a'�>��[g/nt*�R���n��@l<�.��L�s�������q���6��~���E��M��_�L@q�XUY�3���1���+�1yT�CL��v5UO���.��J��d���wi�b#X/o�����Ƭо�d[�dC��"~�d�i��<	�?e�]�U[��6o��Y��ǘ�i���S��}$����e`������|���盓�߹0"ϴi�!�ȭ� �I��&	+��.z`�x=
�Ĳ��P��Z���J���#�Uݥ` ��qT��"�3}��!�w����*@�32�����[���i�+����$��ff���zlg]xo��.(�a�|��uX�:<V{Iz�;S�pj-#�F�l�Ø.VL	�-0Is��'��by�qn ,$�uAZ���'w�m(=�J��%�jz+_�W>�*[��1!M񶗿����ȧ�	����oWڛ�L�=�R���}�I����q�k��́��l��9��Q��d�$�(Yl�8��Op�`����,�����g�IbӫR/��M)5���@�����-Nt�<��Q��+�Wc؅�M��@�(����[��Tӛt��o�Ֆ��5��M�rޜY�#kRHZ{Yڿ_�X�C����|��(�5'�_@�(��~��2��^�nDv�-��~�!��NSh�R�/���X{-��+Qݘ�C��O��N�!JD\��֟�����es���S��� ��ȇ֭H9��&,�h����~;�^J�%�-����G$@2����e%tԀ�NKC��L���jqZ�F(ک�}��5*�浛��"�t㈍1��
ϫ�e��G�|<��ƨ�h��\�W`G�d=C.�܄5�BDs���!#�ذ���o�Ź&�1@�������4T��gm!�B�`�A�ϋ�|�&E��<~
���ת2�5t�4m^�+v샻�>�e�c��.���3�k��- ?��$o���J~Еn�Q����c"��?2shD!^�J+AJ���%! �x=�� ��
�"�.�o5�U�2՚Q���m8[�	ei6�𮮜zI$&�BIb`]����.ʶqp p�Ƿq�{�Qօ��f�y��ٓ�h������_��g۔Fw���Y�����ʣh�̀e�ǭ���+x��U�9LL,���ѝ�5���iC�!��r�-��\���C�0��Z�C��3��;���������ѻ�+�.�'z��CN!&���[�
�[�17�t[�/�&J����7b:18��4��^(��[A���:�QX��6*�ߘ��Gc��G쌡m���'����J3��r���F%N�w��C�\J#�Np_�m������M�܌�p�i�܅��nM�n�ͳ�	,f���<�y�'��N��)��of;�:�	6�"�U�����Q�����|�D�����X2�@��D�~a�|H!�Д�v�&�u�K�|[�q*�s	D��9�����-��������WO�Yu&�-ϯ�i��-ߺl��`0����D@vh˷�� ��0�b�ɘ=���٤��(G$e�S1����\�+��s�d��6KظU��c��*���.�49\�eu��-�ީ�Tv8��Y��)O�Rw@Al;��/|felی�6밪��W]Ւ?�n��vN����4j�!�b����w��c&rlaPN�f��b��]/����*�yB������ޒ��H�4����{�ɼܓ���ZT`�q�_'v�w$��灃LO�#��t����z�̕j�!�n�Į����f;ᖠf4?�?QS���\ȑ��\<UЏ���4�&��Ix��m�k��jl?Y��������vt�[�ƽ���%����Ҩ+g��~���,�G�;�x�����$t����B�I����z]�UaQ�V!E�j�#3�Ij���ƈV����ֲ(]$.q�Z���#Y���S0�t��ax9� U'��E�D)�.u�z��[C�>q"��A��/e�ά����5���Z�D��}�Y��{��{��$?4W���>k�a���dd�._�w�e�PY��^7����)�-�|PX��b�������	�'2����$섣5�d�d� ~�@UN�%U�4p���dk��)�n}�Q!�Xg�R#{7��4]:��ql�����u�"��)�M3WY�I��,�ǐ���Aa�1��+׾���k�P+�mz���u ?ty���]����f����)��MU�����L�}j�ԟ�C��NAz�p�Om��5�|��U�4��sӈ�,�3�,L2�Nv�կ�'�48x�K5�����#m�Ҁ�:�pY��=����P������}����T����~l�e������bF�g lc���';T� 4V!��0��,+��+8̶��ϿU�#
ezX��K��69� f �5���k���B^q�Y�-�0�erfA��E�_v���>�Q+n�
��p��1\�mF��>���ᙈu��^�LL���A�������B4ԘB��ޅTJ
��ۿ�i��-˶�1��;4���\��	z���&��W����H��;�u�G/��� �T6VAeA���l�Ϗ�s����K<�~�$��ڥ4�Um0�+;u��{�Tk3�^�B����ܗ߃V���5Θ]%Mjg�����㔲�*:(���$'1m]��(b�({��p]����?�Ѕ���?F�$�<���=Y=W�E���y˜�Ko�N�̎1��퀗�)�z��e�8�@������iUCO���q�sh��F����vN�mC�gC28�������<�У�`=볛A�+�m�d$���#�#-M��7�*�Ņ��^`��6�(�C�'# W�5U�@�[Ŕ闞��q�k� �pX�Z�8;וЬ����<U�-gr�6�uD�$)�I(�$<"�ȋ���L {-�_��3�"\��D�$a�r��9@�篕!_�,S�*�}{ ��=�z�h�9�r��3�����sIJ\�����u��h�w*
�A���j���L�A���GB�B⡵��˝S��R8���Al
�%
-�0UWH�p}i�𳅥 �*�u�*�v�eG���ܜ��@ܘ�Z֠�V:m���0�L��;w���@��=��n���K���l�@^>CNN��4>���@K42�[4��|t�K�sְ%eG4T����L8��39�Di��d���Kh�Sy�N��[s��&���O��2(8�[��gQ���-Fh�ABKZhf6��F�&<8���<���p�bG���I��� ��1�30IX�b�TnY�h�G�?d+�D[~j��ǚ.���� 
IMvg�K�lط�Nx�F�^9v�nuܒ��![�m3V�H�2q�݌���ۣ@�0(�.��3��������Pt�xz�����N�Zzv�=�Q���
��&��M���Zk��Ք�S�C���Mϩ�� 䕘����=w��E��3�5P��P�jD��v���R��Aq�_n:@oq�Ʌ"$��Ӌ�#�A�+x�f�*#3�vG����q��c�uK�w����`�Es����s���r(U�kR�t�_&�Q�N�(OD� O��8�-�6�O�WB�;��vo��U���u���IEK}]�x;��P^J��?)�?�ֈ{��|�|1*`�s���͑t��Kڶ�]�Q���h�O
XQ0�
h�#A	�7ȉ( ��"��<���M�<�0��׶���L	I��H�_��e�Z=��&�@W���Wu^P.N��l3�ǌM��Nv"�G�=�#�&�����ge�`�`�]AC�h3����B�a��7v55[���qX�\&VE�@|��9)A�f�W��	���SQ�4G�_��bCõX�:$VR�u��g�!(l|q�*l���j�ln����h��7��E���'��d�E���e�;,�ޛ>i&�*'d�M�4���"v��4Dd�էX0?@!RV6�xp�Z2%��<����4L���p����ū=�)}c�ێ}/���豆�X���Y��V�DJ�8�W���*	����,��$Lh�������_MOH_��6%���*�o�/��KGI��\(�U�ZU,;-V���)t�{�	xO�~7ʼ=����1�_�7f��F{���;��~���m�OH�B��˟�G�P��8'
.Q�~(.2|�~�v_V� -�M)�yW}�>K��n�PA�y�P�&��S<�2��i.O��H�G��0.�	0J}Qy-8ϭ���s��_��'���m�Mc/=B�6+3��|2)zk(�}�oTxK������������c�;�/�:�qq�acb����짓�n���0oR/*��`+X5[*�X<���
�/�����K��2dl}���ǆ2�R�SY��7~9����>�(T�]��;	��,�����_������1��j��v�Zj��ni�Y����Z�%N!���#n�i����_,?$E���*�`ЋC���ޙ�:�5�1.�H0��G˲�o��OY��>�� �-��\�՚�����L���'�P�Nj��+5gf1~�5���>vO��,*�7:�~���[�����O�,V(��37+į����T�ٝ��u�5�HD�0�V��(�c�j��ib�e*����R5?P�p�1+w�����e+���d��֫$����͕�W��ܒ�'J�O��[	M@��i����$>�2��8ޥA����E8� �ig�ל�@r;���k7Df�	I���خ0q�?#�^��v8�s(��������i�;ϰ���e+��U�7㊗p�����P�������09]'8��<��5VFxы��.6�4��ʵG,�C~B�(�}#��<I�?$`�^��@�&�o�H�����aX:�5�� �)�:��+͍>��`*�Pl0�]�߰���K ��r�-$���hW歘����L���I"ud-̺���~y�g�j�A9�U_�J�uA� j�E��
&P��c��\˸B�e=ͤq�[3�w�Q�a��� ~�>nl 7�0�ETE��9�8rE�^�_ �ۙ��P݇n�Ir��eT�6~u��
����WX�Lŕ��tK� �F��;{������L^H�N��(;&�d�X��;z��C���&��Ξ�sD�{�#����EI�i9��R�VQ�SC��]_���p^iRYn.��_�St��l�A�j��t���0D��'b�m�x��P��3%����&X�O�	�~�жz΍�ρ?	��m�"�z��������t��!�*8��?d5���Kx�E�Y�n��fr3�mx4��S�A=:URm�FwQ,�U�	G1Vfک��%8X���Kf�r���2�8L�l��d�q�jW���PPZ��>�Y�W@��/`x�;Is�����b��b��ؒ�*on<tԥ�vl��M� giR�\���U#��g3���'�3�.�;&���o��c�~zkBb�1�ڣbWB��/�;wʍ����mxo����F-0��Sr[��'���sFO� ��a�O2��� �ta��_V.?|�rG@x�`=U`M�"~���zf8�#>����xFK_�K����k�m�5{�y�����<Գ�Hu��}�����+��0������Cv^��r�z�\��W��7� ��^�<tV�`?�nBv�y�ƕ$i;�4j;H��ǣh9��cǩZ+�j�z�s��͡;�a��C���(i/��p��>�ٛ{����;U��O�I�jj���jB��YH��	� ��;�@_��Z�4�#sJ�|�p�UC�w
E���ە ��͸",� �w8�x
<CS�>��w3Ym�Q~d���(^nsj����{��m��U�o����?����E�H��ʌ��늽�$�R�g��a�������!�g8nG��&�{v��;�dT�O�*�L�y��u����?�զ������&��#�)��H?|��J��CI�����^~�nC�覟��ܐ/�b	���?�eʍ�p�Cp0�ˉ�>7]�5�ό�g[=�e������m7|��<�a^����0Z5�V�ϸEW<�T�N�!J�y��'_����G�]��%誾$����"|ϑ���<��)�a���8�M7�2��sQɞ�R��<�^ ��v}.i�-/��l�ym�5���_���I��W�-L�|�O���c�+2Y,q^��R�)X�,q�Zpo3�a��j���W��ihO�5��퉂�v�b|���_b���)�tS����>����2b�D�n(�y�d-������%��G�g),�挽�2����<m�ܵA%լ�T?ꖨx�L�� ��`�Q�`�ȼ���cPdkP�-&;M�斷H���
�_<�K�<��{���R*_f�B�<3,���?�n���ϋ��w6j��*��65����T��p�~J,���)pQ	%
�؝_m��!1��z��MJ�+4��b9��~&�x���$�qi��r�\<Đ,.�GwN�0�.���.��Q��#N�zV&Q�3�t��LT}B��[ �B���t�r�A3����8�"6�i��D�K��X:'9=�bTП����Ʒ�gD׎�5�|��ԏ<�%kE`������9Rjɢ��ס��'�{���٧Yfԯm��F�f�Gw�+v(Y�����7�걅�ڙ:�|���qD�n= H��Z!�1�L�ז�e0��I8��{6�����2sQ��*�}6]"�# J���Fe[��4�6b0������z��H�u��(P��4���œ�������{j*w_�u��v���{��9#n���9>��W��A�xg3��j9K_����,���#��Pi�b��6|���4��u���:N����oj_���t���
�nE!�Ǆm65�ۻ��J��ݘm&��'NH�,��CaS ���|��fξ�8
	HC��|�/ÿ,m��#��`Țl8��m��%�x0DK�e�XPH�1"<xv�Zc}w]Mm��YU�~J�>���7OE��r�,j@"~���X#�)}��y�$A���y2P��r�[�x�+I�)�h����;J���U3> xd��{u�-��??^lx6��9��}����Oq"Ɂ<qŀP���U
G��R��;����z�򉓀�Gؤ��Q��L-�����=����SM�9E�I
Xr�I��K��O����nc��~~5i�\m����GC��͒����v�?L`{>�H;��cca��c1�12�̈́{;`�Uf�n��N֥�%|��@V��K��Biac�	�(�K�QSV�>ܷ-{g$rܗ�������\��8���j��?���\^��Q�ڣ�}�ٕS5Ab:s�#�b��Y�sw��D����[�y-���u����A<):�� �J���Bf�����Fj$�[�B��@9�ykÕݏo|�������?r�^��!x�P� /��r�M&�i1�4�|�{�&�뿕3��\�>�M�a�sDx{:>����b�� �ŵbʥ��D��(����^S��W`�h0W�?�ňv��$A88��b���n��;�V,�6p9����D��hG�@2/�t��_w�T��z*N� �����7�\����0���İ�- ��07�F8�@+��JAM�5����_ť ��㴈FHc#�G(�p�>��	q$>�YN&P�稞����,�%��7V�P��_����l[�WI:�{L%��(#��n���2�.ܤ�nj%���M�c�d!���ca���0�b�+2� <ޜ�ۭ��AT��zwDg,���}�2X/`:*����Ϯ�3��%W\�I��*M�7v��Ǉ��\�2��;��<�L[���b��Q;HmM��a	�J�����4iQ����gU�%���1_Meɞ�	"-�,[����z�1 k�Ӥ��6����W��D��(�����i���8���I�7�̒p���W�e���R��:�P����,��t��2�&Cn ���jM-Ά��yY6�I��N��BM�B��&>3zN�#�}�|����E�Ph�k�+��^i�b70FMݾ3�an��g��5]��U�u�u����C�d�$I�.��p6 J�W���K(�J�-���r��BR�����sg�Q)�2uL�gM��s�⺬�jG[�9Ԭ���Rnҫx�iEh��=F����Ďݖ89ݦ��9`�(�*F��۴QE������\=���"�Y��nQKDJ�!�)�~�ty@���h��D��V���P~���
��� +����+��cuI�B�ݧdƬ]�[����~[�l��:H��M��pv�.b��N̫�)㥰;����zAY�&N�{�Wy�^Bw��B�j7���E����a���}�8�OG����j�c�A3��a���m����������Z��!�-�R@�M,������=���x"�l,{�s%�#���%����,o�{>\�ʚ[�\���<g�p%��)�
�5���.e;I[e�kh*Wc+ ���NS1���ި����@���֨�C}�g�[��)��i^�0�Nn
���<���SBB�d~��¹��x�m��|2����%zM���訆>� ݜ>�,����Ą���P�j�@��)q��X���RD�'�п�]��]f�#똸2<^����V�;}0���'e����Rߤ� Ƚ��4:@r��At�`��~S��hdS�Ǽ�5}��ĳ �;�$���a�ֲC��,� "%��� <K�PTF��Y�}��E>O��ۋ�~n�W\1(q���8qi�L��Mu���������Z��u⌔r��=�&�&Wq����H�`��Y
�wYzGou�|]�3�6L����-��i�Q�����i7���T��'�*�Ĥ� ��4�W�6��+�)���x�cY��2���=�C;��c�)ԣ'�#3J����ЫN_��hX�U���5���Q.	ٚEEw�O�B�w"ʉ¸D_yԞV��f5���=�Q��6��x���p(�d�c+�u����5���� .���i]r����ԥ��^�|<�X��!|����Aa-��5��M�#TP�R�����+~˅�'g������r5������Z�-k��.|N4������M�� �xM�����-�i����*��6@9�7Ղ�gS���I=*8M�&(��	T�2ٹ�?��c�� GTϝ�T�A&��֙����F^<���`�n�#^=(Џ2^��)�w���_D�3w�-�x��c��mt,yq��K�2w7�2yf(}�ˑ�T�L�g���Rcs\�4W�isU�U��u_Mo����JN)�x�P��I�ɤ[��rb�*�K;���-[��^1���M������d{�^����k9]�h`Q9<��rdF�����ߚ�1Ŋ�%�G��0�͇�b�t#ư3pW�2����w�B"g�6I;��uNn����������0���[-��n/�F8�<�ɋ��qƿ���ub�ڷ��J1K������x��N�B�;W�����S�Nv�Jq�@�v� �V�ϧp��£C�z5zeHZ�sU���Е�_Lx�-;s󠬖>��OdC��|�>$A&%�w��N����'�=��><��2��	}���s��;�1�0q�Q砃�Bo�4z�ކ@�4@F���N<3�,s���X���7
ڶ��2�����/�1x�v�"PS,8���B��4^1Uf����;qش��_<@k<�fDd�� ���yc����ݏ��>I�;�ǯ�H��t��l������b-�ډ�������������莋�g�S��y���Tբ��T�Β7NAD=bJ���˙C�~���"�9�����Y�D����;��i0�4U3!��K��[ӝ;�P��3f}ћ�,��u��R�z��aF1��ѭ��v���M�}�}g��z�>cΜ�wF����~��GR��}qW_y��ڏ�/�d�ymV�eC�_�� ��q��T\�Whlܩ5ȇ�<�i2��p��XV����g`U���|X��_�����+}h�q�t��i���[S ��5��1?�}
xW�L�ŀ_�P��@���p�w؃d�L���Y�blfJg�?Ɣ:���]����� GJ����^ڰl�Y�V��s�����sH���x�Eܭ����}����
!(�D1荍Bs�^
K�E�W����j4]獛vV1 ��5K�J"}/��=�*�@�בۍw�t�/�<yy� zL�;�ѼzUA�IK5��.�C�4��x;��R)w�zm^����'N?�}b%Ъ��K�G�<�`��q�¢c���fm���A]��C<�+��1#�콴;(6�C��]�^�*�1I �2+]�?{��v�'����zB��&0"q�2���v��=}�ٵ0�^C�t����ـ@��t�m���>�$"/�ڎ��L�e�������9Y��H*�rK£��XY`LS�<���Oru��w�١��+��&Ǒ��3K!?ǅH��D����;3��T��7Ϳh�B[J�׋`a�����%~��P���Q
S��#D|�����4����S��U����;��!��n�>t��!5����ë��P��? Bӡd	������4�� ��4��ˁxq�OX ��I�>Hľs�LD�ݝTɣx���l�ؚ���X�(���̞�9U6�l���`�j��q#�@F{>Vp
/j#�6��4!�|.��x��'�퓜�(�I�1�wL���eBʯ� Gm�\g��.Tw��i����c�@��x�o��~���Y_�,r���P=o��N��f��-�d/f��u��v�$yu����Be��T��GB�Z���� �vh���ծyt��3�7W5z;0�vA?!NIc�h���W�>�V�x��*D���\�<�)� ��e�ժ �dG(Pj�%��HT�hn�1=��1�%3#��&��3-b��}P��xK�`*J6�i� �f^⎢��2}�V��Ȥ?8C@d�������UƑu[�*$Z�YL�������Q�i��m��zmO���l91�L5��`����9K 2I$�WLy{�<}��E��dԓ�B�>mǇ/���]f����c��2ǿ�H�ш2M~'
�¡�$MNa�e(hl:��佛�� �q'�ٖ�S,�;
CY+V;�f\���s�t2���Հ����$¶$G��ۑ�]V���hԊ��a�� ���T���4+���,���Lӕ
��$Ȱ����y�
���g��x/��<����~j���:�n��U�O��ʡ�����bלL�۹�����siI���[q�7F��H�ν����S�M(����:�
�U ��-l�͇b��(���f�d�}��+ac\��L���
����l��?�b  �w^q�v����l�_���ƀ�,Ή�����x��6��8�o~�o�2��H�	���O�5�P�a�"m�X�v7�0=8�Mw��4��÷6���AP	�3"P� 
J��L����2"�K����&	�!p�1 	�?I@]i�mVن(т�o��p�` � ���$$A,~�@-�%/����Ji̑��q����\t���2���^�s<�2
����P���h����8PR�ϲe��i��H>�<�������4ǉTn����k�]�D	}m�M>(����Ef�*���'�{��d���A-+[���Q��ʷ˱C��vy���;�O�LN���V2�����P�!���\^{��Xv�CŻ�s���⎦j�bѪ��B0�H�g���<�G�.l�n�W��hb�bu�'�z���\���o�~�.=_���z��� ��|r
�k���v����hs���F��p6��k���1�PG�[���Z��q"��T�#bq3���d��ƒk?d^ħ�?��H�'��s���F�����n�Z���1TF��NP;Y4�����\���Ҷ������6���a��Γ�<'D�����[V3�,uۖ�$�Z�e�ƨ��:
���a����S�5�i5�=sZ�~h~�ͻ�t!l�8����mx�)Y2��U$�
��֜��ׅN8Q��d�4��]���x�N�����ANx%h�Y����$��7չ/��j�_��$y�1N�g��6/{%g�Ǥ��F�~��d�g0P��	�w}Pd��U

�\c�*�c8��J!cl��rT���/��I�ڳZ���O�[����l9j'/+�>�ɡ�.h�@ٔy���oz{V? �9��\XS�34Cj���e��C�#a�A�z��QA��P�˴�m�i70�B��R+�	�ՙ#XVxg���B�-߅��xY2ZW��O���L;M^Ia�d)�L���� h�5#�r�"��C�Ϭ��i���Z�l� �IW�=Ԇn�	c��N~J[�3� �+������ޗa��/�F�w�m���=��DpL����a���E_(E-�HP}�m��}�iY\�n�Ӊrd���ł��9���֦�M7V6�r�S�,�o�㓀Nc@N�e�<o
��o%�x���撕wG�
�H&�����-�&�}��L�\u�(-8�� E��:�_Au��P�܅�C���i��g�|�����X�+T�p���`_�I��5�ai�c)�n�=a��N��'5;nhk�_z�Gw��n�k4ϘBӘ�Fnkˑ90X��׏	�=�S�c�}�4釕�;�d�4B�{p�=����3swb��~dM���[�x�Ы��^<Bsr��v�7{"���HZ��%9/��GN����}5�,��gO����^J���WH���ឈ�����{�1��V��M�V���,�[8��lJe�����O�x/��	O~���D��?�� G��0M�0?ݬ�9cs��i����𗬆�@#h�>Ţ%&���r�]=���KLcn�0cV��<��j�߲+8�� Z�
����.C�kY R��̟u�<��b��2�A��*d�� ��EjE�i?���������n�VN�H��4�MR���*�3������
&BV"����5X�#`�&,�u1O�K��KT��Kw�3w+d$Dճ^*tQT��=N��N�òt%�}V#��������;�t�;���M���\c��]���s�#���f��w�"�M�ڼ#t�o�͖OZDP�C1�����d�#�
���3m���ʴ��M�|��C!��-��a(t$��@'���uL�H��/*+��C7F
�Ӆ:�x�����n��5�jh���-%��l�!�uj�ш��Y,'��t:^�̰����� ��*!I����x�]k*�ӑ�Uab5�L��ݷU�u��<�4�?�M��������"=��ϩE¸�t��I�y����$��!�2��C�cae�����kl�|�&�Ӽ|j���Ρ ��kO�n������Ū�����<髟�HG��&�*m�b:�?!_|�່��h��.��-�[L��)9��1ej!Cp��
�������������|mP�y�Rw�ad�M�m"T���*!Dl9P?��a6]�y��V]\;�;�E��O,����끂�F���(�f"�\^��vp����I��)|�+��6���A.�W\m^U����a�&��Np_%��,�2��Q�	��_�榜1�jGہtubgF��l�J/����|����U�k�U��B�v������K:�'���R:�Dp\��֍]ܲ#��s��L��p�n`����R���$KF��0�'&J�>���F������u\�H"~/m4�ɒ�(/�ϡ&s6�L��ƃ��>����Ғ`i'j�2���XKk���(?04�E����!����E��OWcN�뒂��q9�딳�U�%� ���{�P��m��l�b�G��f\^K>^Nx���� e���~f���A�|7�����R=�82������(qG���\�#��i����Cl�E����η���H��fSa����Fb��\\�J�1�OfV����6�yo�����f�gb��?z�U�U�R*2�8a���M�ǭ[ܷ>�c���Rf� Ύq�-��sT�R�	T����;`Ҹl��E��-D�N���6fo3�
����!ր/g�h��q��&�_��ty��(��BA��J���zB�Ŵ��Q�B����3���T53�����T�%��=�];,\� ��]���cP{/XW~|��lܘo#L���SvP�gj�׵ʼ� i�y�V}�9/\�����y�En�K�9@���J���6�h}�"j��/Wcn�!�e*��ٙ���/g��)%�_�%��`-��=�ῢ�j�� >��AX> uYY`㑇ŷW���n7�ۈ�G��N�x�ou��f��54�hU��w�h��B���ẃ!Ӳ�}anӎ-�O~ܱ�\��ُ���c�Ŏ~Qa ���n=(��{�4ATIgE�N��L�t��
�����*5��RjȜ.{,~?�s;&�NS�H�����QD
��ʢc4�uDgd�5��е�����$�jj�������$��c��I����X���`��X����3�7�V��=H����fz�3��?O��-?s���x9��x�9p�b�Fo�n/-C	/���!0��*�{��x�R�c���#v����Y�bY��Fg�ArL�S5��Q�G�xU7GB�RO>vQP�#�{�y�wI0��D:�V�Ef=��pJx�����ܧ�_Q�M�Mۍ��j=� �G��̪}X�U� 9��nV����R�r
6���C�k��e?�z��`��$�83w|�K�!�`8M��vfn<黰� u��#z�/2�|��h��5�"]S^a���\o�|�#��@�
�h%����u¾l�.��+�}�Iy�ubU�P=K����K�(���"���p-�(�
)�fI�ä.�hd�d�b����� ��*ǕE�cD<�'u��\��l��f�znP!��	)\��U�X��2Mf��1�*B�S�
��#(_nb���,�f��c�Rf%��GE�
^wI�ec2zGL�#k�]ED��wRɐ)�o�)�l#�<�'��w��d����}��7Y/�t?5���hۏ�>֊�O\c*�CT�(y�H��xVY�{*�,d�H�\��y�szB.��<���Z����ј���Ee�C0��p�1�xN�m�q�S�� �:��g���:��5&�PD�i����dC��"�g �L#X���lf�2d��Vv��9���D4�̐��@�lw��s۽���.���
.�}���/
w0T�'U{]������^YH]�tos�fL ���S�~����Q��7��ꏙ��iK6���|�A��WH��`eW=\	��
��/Ԡ��Qdjb1�}�v���;�ʦ{�3���+N��O>2�/=�õ�߬\ӿ-���eL��b>��?�|��џ�3�yކ`'� �%��q���y��U���<PW�&
�6�O��Tr���0�j�>\�GD�ҁ�"�0[ٿ�ם�Go8��2_vP�/z�Z�kC����"b��'�[���4RAq�]���Md��-����̶�0���YƧoo1׽��!;��'Q]���t"au����r@�4��%�,F�I��@|���ܵI�g��k�%dr�ao�.��8�������8p%^������f��s�w�V��� _�v*{C�a2����3�jB'Q"��I�����N��N�agy/�%�Lw�\�}��-��e<0�4r���@0�ؑ�
c��g�,cot�<�Y��C ��crG��Y�_��X���ş�CMJ`	W�ͅ�`i��TK讕��9-PO_��d��?�b+�Co�Q�j�0A�H�i�
x�չ�?�A>)������n��\əac9"��Gii��i�!�"U^U�<[�װX���I�T(���ޢSY��ظ�̢-�G�Hׯ�W�Q�����`�l���vg/� ����* ���D�f	2ZG���5�h��1��5}�׭���B�=���ő"�;x_��.,s9�)�X��ȿ��F�dW�E�%pl�#�wl߃)��mY�������,���M�����Q�|>;I��P��e ��SW�6� �4~l�@���jEw�GJ���?���s��&q��M�у�q!��1�XB*u�-���l�1��,@���X�Y���N�	iiS��0�7`l�jX��7y"�I�g;�� �q� $�'A�"g�~�4B[�3��3��/T�2O�I�J�o��`3@����"s���=��tJ�f@x�M(�)��>��݃�(�2�2����l@)v�Yd�A��Z��f܈�♇0���;��JU	��W������f8\Lt6>U�'�ɴ:ś����!�)�B�v��L�Pqj�t������(J��s5q��Rl�N#ҿy|cB�"�Q��$#tt�����y����	�-�S�B�~�:kb��c��Ǽe����\�Ok���S�6?h3�3u[��!�6U,�'�az�ȝ�Ҩ!,��K}��*9����~�Pn�V��p�3�lЊ#�4fr�7�R�@mk���rxV׾�8��͕3������ff�H�Z��G �u�H&��E��BԀ�V���A�V��������~�+'n&��3Y�kHe�"�b�V�6X2�iEG� �@i
c{����z<��<�a��Ιp�S�C*�mH�רF��_FW��;��.�P9^QI��w�aԌ��J�`Xy�p��8B��Ԉ�r�kF>e�`�a��� �����pÅ��$�Q���eG �ئB{�rT:
5(�!��<��P#���A�ή8SȗS?������i�U=�Kx��� ܌�o��1tL?p�Q*¦,�t��t,����c@��
�a�κ�*bJ��h5S62��Y(����B�?]�AA�Q�8ʈD/"j�a�C����ȪH�q�"=L�xZ�u�*����&�?��'g
gz���&,�{~��`�X��q��ay��ąi-C�&��l�ݟM�DI=(�"�Iy
%dC榆�ε��#��n������~d1?g����柞��.R+�*�<��=��ʻM�EN�l;�clKe���f��*�J�2ǦKm�ޔ�C�xs�ہ����g��\�ϋђ�<�i��Y�t��~)M�cQ�F5�����ƞD�4�^z_=�@>��t���!���8x�v�h:�X�~W����[�G�M�rk	F���2qx{e�=�s�)�O=|l+)���z ��E�E�_������lδ?~JȶgW�N�h�Z�J�q��p{�H|��.�K΅Q��Ų�C�e�o�v� ��]���~���b�?��Ꮩ�#^,��p�܆�\��@�Y�?i��_Y5%6inpT�.��\�7�ѳ��~�æL�Q��qL�{�_6�o��4.!�h[�|�;H�* �p"+��S�렖�d��,_f�)4K�+��S�]WLl�I1*? is�3�����1��=�W��y�c��P�������!�8�	W��7����X`_@�8���UfG�Ztys���7ډax�IZJ='&ܮOH��uv�{H�e��� q�3��`���N�{��O��I2@G��e�/]R�G��r�0Β���z����)A̡&ҥ�KzZ������"� ��[�9���3=R�g�]�<��"w�jR��B�A7T�:�U�6����})�:��^a�vFȀ��x�lַޒ��z�' 7ǀ��z>��V�t�Z������P�Z��Kz�(U͹��Wf��9h���c,CC���	b���lm����0�B����Hy
�i�����g�sl�d��bڸ�`OE_�S<��g$�o�M�\Y����&5�c+0�K>l�M��ӷso ����Xؕ�����Վ�  r)//�~��ie3�esY��t;�f f��|��;^BrR��˝�[��i�h�J~3r?1�u�������B?<?�
����6L��yO�]i]~����'R�_�I�/A4
�5��I�3MxE�Y�W�*���Lt�8i���x�
��B�?,#Vmz�e(�xm#N]�l R�
F��1EQ�A��\EG5��U�l�šd!+_����ʢ��*�I	F���<2�6�?���dm�3��^!��8�����Ds�P�ю��W�9�dh���J�Ӎ8�:D���a}�~6�5�0d�|�o� �-[��^�~	���/�ݷ�j�����T����|,�j�69�[9!r�,�4�Õ�\�ihR<�Ǵ��H��(=�Q�⨣��qH������������%Z�̷o3�[��k:�kr�P���:�Q���*�o�����U�&��M蠷Z�]`��PM�r��or�+�
{�*�g�뗶_;C�!�X@��C���r�Y�$�����o�M�����X^^�q�Ȏ/,s#��G��׵0	T�ҳ��fH��EZR��f	���}��)�՘Pa�Y;$�B �;jiw��/��c�@��s��ܤ����Tn{�?Ӣ�NYQ���Ϳ�Sn݅y5��Gt:[h���#}�IQ��{���$��zY��c�z���A�x>O��WjU5^ �d�3?Y�d��ckW��~t����_f�k�u��=Q
�[��N��������S�zm�}�n��%�S�8�@u��8	�|l��������,��TJ�x����� ������~�ő9���T�U=YA���lb>���3;�R����f�J��-=��2U��c^p^�ٜ�{��!w������*=�u�i#���(s�규���ßo�������W:�!�����"VN�fA_8�3�:��ٻ��g���w�/h���<\#)��4�8ςcE@��r�땪2�{!�1QF߉��1Ӱ8�T���o��i�*�B	������޿"�X�yE|Yǘ�G�?��"P�V˔K�A̬y�c���e dw��������XB ��d�}�b��J������c#ronF�i�@��Ԛ�H��1HОLVO�
� <�A����`��S���]F�{��.
"�nK�v=6V&VD���rD�!�F<re��M5<�N�I��	�F<�#���#%!�_r�A���7�(�r�j�}��Ŏ����Y+�6�mǒ��x�p� L�v��m�Fx�>s�Ũ�B ���6�r���l���/�ȸ+�G8}%��`�=uB��B�OQ/ �O���K� �ĩ�G���q����z�{2�����%�m�e	�����n�>! �?*�_тF lK�N%#k�����(_s��T���n=U%��)e�e%xsY�Q��X9�	�� A#�QX��sw�����o���ǖB }�I������yK��%�ɕ�3D�x���zG��Ωx�
�@ b���6�&���(�χ�p���%�- _7	��[İqb��u��i5�vE�
rV,΀��A\��p�mHzP��qR����8_l XMO�Q�O����'�UH�;}�R�>��o�ϱ&��� �Uӽ5)�J',s�+�?@
'�I2��k���L= #Ji�'�Άo�1U)�=�ގ	l�O_���bo�����pR��97}<r�XC�4M���ј���b'����s,�� �l�<�R+B�jF��T���8e�duA��#��>U�ص?��Gh��C8�ɖ���O�D�LA�9c���(qS�ɤ矂u�̧V̗c���Nr��tÌ$��Ѵ�P�g�'�x���P��S�!�s�I�r��l���F�΢��s��)���#���%�c�!�_��Qm(�+�E��UJ����qlH-�8;�L��DS�FBҪ9>�S2*��m&\�@�v�m�Y�φ��1'�Y'L7������,Z�>�ęsw&����}��Е���A�������"��n��t[G�{��p�ʽKB(�w:|���w�]�����Vr C���H�+�H-�j���mHV�����-��N4�o4���a�է�A?^g���* ��É}��ƨ��Z��;��V�ק�����y�p����no � ��K����m++Y��51mL�%(�z��b,]��!�]`*��[T���*O�ӏ9<�A��qw���h�Z���4�y�@Bô���7��{�*��Nm�I �9E������þ��oB'�#6xD���6Pa��e?ܩí�����G�*ݾX�:W��Ձ���s!� �dj2�x��z��Ȟ��M"1�?�ȱ�W1	Nq9���[�^����k<_S�$n�H��bKY)Ân�D͡�qbn��Ѭ����8mB��7���o�v0�����Y���T9�*P}R��
�����_�^U�3ua���j��ʑލd�-���e�UHn��my}:� ��)�-S�~�L�1�0T�i�M��jz�j a�Ը�T2(�Aig���)�A^$�ҥ0w�~(?Be�������T34�@q_0�*����N��>��q�y�	�[��ab�.��(����r^,i�Ő���,I2_�uZ1za��n$�ô��A�19 ~.O�����iM��_�L(�k��H���Q��Ez�����+�V�--�@�gyqp~���<6�4f�N�������A���Yx���P���aY
�6���8��~��y�in}Yp_�m��[�o+�u J�2o1½�w�3���΍��@���E�*��I���y��1�a"]Ʉ����6uN}a�([i��2cuߺs�S��/%M�z�D�s���C�)(���π�J�8�To���x?v�Q~�oH2X����]PS$��E��n���}J۽Wj��u\�Y����2�^6%/�i/�e�=E𦲌G�	Gi�յ��U�;t�_VN;�"A�d#�2���G��`@�X�lh5M&У�n*�R��n?��.��,�],�N�b�:?�mšj׸҉o�»��&AM����p;Qj�q+�t�@��"Oh�c���_`��*���t1b
[ϊQ^��'�D�7��νmj2&8|�S@G�\U�Ѣ����'m���8�����w,|ZJ�콈Rm�7V�CU�G�5&�ӣ@z���uj�i�(bW/V,����ZLdVa.�d��]�k����!�qk(7H9�Gt�kjA畣Ȩ��*f���s%	�
ҩ�i@�e��h���$�ՏхQ'�%����.*��1��G[���v^jxҽt[[���q�xQ���ꗰ4�88��A[Z�zPU�n�^������{elj��\m�M�&�poRl��l�\Mr�=T���`#��o� �vY�����x+p:����������)��xF:"��5F��UD��i����w�(T(��A�{IgNHD�����$:V��J/$*�T�Y�{<���<mN�'�"��H���|��+b)P1��i�f����[�@Bs~�	 �5O�V`�	�
�+�K*�f"N<�KPk{�kJJ�A�A)c�i�+��$��cΫ�SU-ɝ�ؖ͝
���/� ���i~K��28GJ;�b:��X\ƚ-����9�e��Yf����=��i����#�!s�4��T\��?�P�K�%�A���Qk4����?��/|��@��6/X�\�a+ �Y|xT=�v���@PO����!&;���ٰ�*�@C{�6����Z%I�oF�;�A��
�*t��d(��RO^���g'Y^a�~��E��SP�n���@M3�G�����x�f�aE I	�3~>@DH*�M�u���,�.ё�`e���#Ԥ�����ښC)�Ղ*�`Jo�� ��.c@��\�}QZg>�!���]��h��q:�C2�g�6���#~,�E�<�A�OUh�����(wS-�"�o��%:�����>GYrxg��6��Ӓ++��r��g^���b� �H���F�ٕ�_��>+��P7W���,i���h�s2\s`�"{Kt�f��$z�J�7��)�	�*Ý�H��@��#�l�N���P/���q���������âwe d�G0��65���j'i�͉�f���:����cL������5$����ԅ0�0d)UAl�ޭJ%��z~B�c�߲��}BfY0�}F����������0�}��[�X��J�E��݉�#⽌��se_��ѯ�!��"Ԧh�Γ�f^ɫ���_NY�QU����G�M����nf5o=���ˡ��C��U@P�L� �\G~�����:v�^S"|� h�3J���	\�][��SPq�ٓ��'g�2]n�'�&�U�θ���峞���ٻ�]������@�O�0+��I��,����)9�A@���"YCXi8����B��:�)�SK�7�����b�J<��S�AW�O`�+p�[�(�T��UM$��]tT
�3�v�M������p
���"Oޔ����;O�I�1����tQ5r,A�Ϛ[B�EF3�� �,��.pb�S!j���E8�-j���oV �I�+��9�W��?�0��"���YT*c2��Ec���r��M�����|=#U�E=��m,��!T����-2���=5���p*�'l{@aJ���6��JoTQv���h��9�<ś����):"ik�ኁ�6����I-�7i��6�d@��VV�ݝ,{�j��J�;��(
�(�R&�����.�c������f����`�� �LR7���NU����j��e��%��4�������wI[�A�p`����C�I����$��Rƶ�R�-,�R�A[�`H4��|�܎�;�g�)$m��[yi`�툥�$�uK�����
�m��zu�!����A] ��˯2nJ(�6���*Uи�'�8�F��J��s��Pa���uۛ3[���X��)��q��qͮ�������S_� $��b���X�%��r�ɳP)�C1�R�4�
3�Ѧ�%����a�_�Z��E�c�������f8V_|�ACiyi�Q�ǺX�3����sdD�����	���k��R�G��[����1�Q���Kӈ\�փ�rV��g����<-���?l���e�3<*�+xw��r�<��E��и�+�����nl���H�V)������HE�,���Õhߖ����ɦAd?�5��XP�	2�657�Z�S��lb�_���?���-��R��d���E�����cT�~z�y9y��(��F'�!��y��������#�t�Kk�g֛���|�x�rԋ�T�1T�Mu��Q�"��@W�%��M�㹊*JP>ЏZ��P��dƝ3��lX� �y˓,�?�=A���D�v��15�+xaz�}_�wgUq��˷�͞�EL̐d��=��O�l;(z%nJ§�аn]F�4�������2i�V�.Ҋ^�S�����n~u�.(rt�-���Ê�:��'��Pi�^wX?��
�f��)z��N�hou4��[��� ��5����x�+2~�Ҕ�IǝM����ܰ�!VE���R]�8��Gk����o��f�D���6��kf�Z������W'G���s�#�3 [ҹ�  ���$��g�CE�ZA���x滯rv�#r H�؎J���ò?���$'���l���Ф޸��0:{\O��Xe�;�Vx%����F�J�L�
2	�� ��3��a�F��O0��h6`�,hl�@HLඝ�����s��d��'�;��E>����lnS����ҝ=ll�c#WT5+�Lß�����z2��&Myq`r��c�����̅�m*0}��l5N����\C(���=��ڟ��p-�jV;�(N.� �8Yc����s%�[{b|��2��FO��Q������׭0�����~���T�d�b���Gۄ���Y�]2<[iPo奸�@�9��~S��࡛O�9��VE	�|��Ǥ`k_�zE�d���N�'qh���x �[���	$���8{�=C������l8^G	�#jy�X�	�tI!N�ǞOG�N�*�#5p�=1�v�3����yH2-x�_��Q�u�_�g:A ��ж�����T�R���M ��S��Q>i۹i��0��>ښ4Ǚ��θ�q������r�}�lV���]%\�|��?6�����	ׯ��p��JK��9i�o��m;J�����G`9�3^�G��8F��mƃ��tJ
����0�������X;�~ɳ�eȌ�h�+�z�5��4zj!��w��z�>��\ϐ�P������P��2�N��֎aY0*j�S�*�&�ň��e�8��&�+����"�ҵ��t�bZd8�D0�(�ۓ��y{%�ދ��ýG�$ýOf*t��6}"M�1q]�y�!�|\
&����m��xʤj���D'	�7ܿ�O�_~�6�\����b��I�GB7&�$�c�2�fp�D�UX��@�d0�E�~ ʵK��7�Yv�J69/q�c&�a�7�Q1��4�6�G������r/�5�쯔�K�	�d_P�SH�|�Ga ��q�O0Ē����r-�&odZ�����zt��#��VA�$��0
�}3���NЀ%��d��b�� �B���+����P�g�EЉ^�!���ފ�%�ZI���D���g��Ş���nX�
p�?�p��T�jal��2�G��A��xR�}�ʷ������D���F�A�`mw��?h�~J��x2ɽ=���s���Qz�G�Oe�p�Wؗ����M'L�g�������#b�8Ob7��m��{�(IQ�f��8�k0�+��Z2`�G�$����jdб �9�ȹ�K�B��yR/�Q�I�\�OD� s���;	��ay�h&n1
m�)�XVt�P�C��(CO��'o��ݕk��**���wu���s��.��{U��<נ���l ���E�艹�J���L>/0@Zn�Y��q3�rx�;�~���V���x�f��L��H��ވ:�yTD�l"�X��*=B�/���4�9�����q��<�������p���㘾��2�:�r�p�W��9��]�	�Y\莄"��"y�Y��e?A�"��*��;>���KHem��	Z�Ӻ
+*�?�F�+����B
_`����Pei:�a d)4d�yոZ/�D�p�<�'T�
ˬ�~�QO�bI~~����g@��x��ۿ�eV�����N} hsx�4�Hc����7�O���d�O* �Y�D���I��gQF�l�S�x	�C�pPnpǻC�T�wI��r/hSɱ�a���\���N�xKX��x߷��l��ܠa�8����%Ҝ����`8�߃TȈ7$F��M���)���)L��_vZ�۳��KI\�B,,�*���+����F�c�-���ӷr��h�.�i���6+7��c��]�̐;B��n<z��6C��Dm�<��!���❖Dim5����n����4�VN!p2��&���Ը!U��Ҝm��a�7�=��2	����fǿ<��y�m��9��sࣺ;{�QN�׏/������z����c@G�I}=(Hd��23�Sգ|�1���R��`ߔ��V���t�vh��ri��o(��j98��f����w�]�i}�};DdGn��C�/���v��D]���F����E�(�`^r���/lT�-KS�}::�G"��]�-�z7Y}�tf֩��G�h�L4�@���TCpqQ[��E�����Y��/�80�׋�K>J�J|n��N{ŗuҥH�a�J�G���'���Y�"����V�Iv��ٲ<���wj�v�/:�Ag2�8*�]�LrA���F�K�T��
Bt��v}�Kp�F��ۮx�8#H�,�+��NiX֕#�H��فe�UZ��K�8̆�I�d�:b~��$,��q�Ǟ�Pꕀ��H;!����n��Ydib� �ْ�]�x�蟋^#M��J3��?�`V����'�ր�a��G���^/��f1�� *J��*�_�@��i���7�}�s�ŭC��m�����eZjcB��D0wc��h���[�9e�q�A{+Ar(Q��2B��e�3,B�����:2̔h� 'Fem@�LK�,��%<�֝Q)ϦB0��֨{?ש�kpM�=E�Jܐ$e��JF-K�Ӆ�s��k��H {�$d �+>�ˁ,e#̘	�N��%�ׂ�	�*�/q�;���������e�u*��N@ew�۪��j��Y��ї��_h�Ɋ�9W�_�ù�B�Qbs�,>�E�=�BL�?h '�i��]��k/��  �ͻ�y�1K+R�A� ɥTe��ɞ��h)��&��;�Ӷ����h	�٨���jk����f�[.OӓF'�R��HB��ѩW��+��Z��h�S���U��~I�h��HkS
PLc�l����:�Y�(���ٍd������0��}TC�� ˮ�m@��=�'�QJ��ЮhM�R���<q�b1�2�"���G����+�����	c��0
��d���D�
���<�e�����r7��ۮ��R"J��~�JбX�oˍy����c�*��!����U��F@��bH�zs���/�!C����`Y��	��-��D����
���$�V�)�^i�.���%�3~N<�����ԑ��"� �,�i,t�1m@�S7�����$ѩr�0��s6>�hpr,�0'��	
���\�ǧ's�k2MĄ|p�g:({�v��`a�Za�5��-�Db��n��!wZ(^{� ?������W��D��g��&zQvr�T�$}e��K�MK�, b���Т� ��$���i����ʑ�D����{m	���Z��d�rt�s��o��da��ϡ����Hv�k*qc[�.�瑈�S�6w\�ms'?x8�%�@�Yn�h��rGtIhݻ�\01G�c�i�$Ҁ�:5��Ⱦ$�^�xؖ�b6J�������x(meu!����:��=�����R�U����<�_��`uxX}�x9md�����a�!��rpJ��r�]��3���L�s�;�i?s������XY$k:��5�I����İ���7��p���K6�7�Jp�ML�z������:�̸uZm
޾��?�i"�j�!/�+��>����9q3�w��J��]�JK3:�0n+�E�ʰ3��%a��q�V������>�xĤ �r[!���ׂ�z@�
���^R>:�����L�Dk��u�OsG����|K�����;�ڵJ"[f$K��NW����Gڋ%DP����
P�"���A�~߸�@ҁ���
�C�$
j���A�;�-ju���?�����.�-��.b�Ԍ+'��8ȇ�� ����Jm��34�+;���=�(n����533:ޣ�ߪ�Fʘ6O	�{�rN�'� ���=�H��!Gl�OZ�n:����gI�,@��q,�:� 3q����~��mOTC��X�'Dn�J�8�Y���\��Ѷ����ݨDf��r�
��%Xӛ�U��w�|gG�!���nW!�^�N�]�'}���8�K�� �A`ʡ3I���6l�\F�*�h` #�*7*�EjP�?����$P��q��i�q���B*�Y����F8��;������ڳcb}�K����]��)q��tB�9pƯ�_��k�Y&��㙍n�m�^3\6���X��H���4#�|�;�Ąd(W�ǲJ<�v�cm��3J5kX�,n�-�[�'ڑE�(����!����mM+K��q�����<'E[b B�7	�%��* ��}a0p�Vô��6$���t�g=�U��V��g3������3h�'c��6[K�_C��r�9��4�YϓY��
Is�q��G7p5US��Wq�ɺ�r�E��C��@�b��	*�k~�ŹQ�}UY�*�)~Z;3�����._e/;���S7ɫ�	�|4���YF}�Aa���@N<���u ��E��=/������o�R�2�Y� �'�/���)kv�_��Zz� t�����ΘߴvB��q�Q4mY^�.
�y6^�f��L�J!4O�'��Ak���?˼��*����TS酐�A_�C���)��7��sW��:��g��0�|�$��Dbk@��+)��>y����X�[��hĖ(Q�
��m��v>\6�{�k�?��r�TE-��s�)�\���=U3�������T1�C'}8P���l0����/��{
!CwpmE��`�zZ�z���%��f��N<������:�bm7�w-��Gˋ�UV�u�XF��Z��i)���"�+��~V]�Nߦ��ی��:P�
K�N���}$�T[Ӷ�i�eK��
ǆ3��R��^B��B��e�5��]���������>���:)��%z[��K�`Dvl@J0_�^��ָ3��E��}��DO��1����[�B��w�灥��Ы4.<��$A�w0[�1t\�Wחw{�g�2$����Xb�M'E��wJ���C�Xb�����&u�h�� �f�PKT8�tݾ�qJ27S ��K���4��&X�l.�'�[�-a}�!g�o�eQ7�Qa�h����3ox��,�Lѹ�P��X �D�֞�J(����
ˤ��5�q
�r�a�A9����(�ل�)�=0��8dK��	�޾Fp��c�9-jC�(5���������Ħ�V���{�ɽ��{=��k����2P��?�r2Tj�爳����8 ���<jh.�+��|�)�w-@d�ʀ,��4�H���+���B!�0�B?�n����B%��E5"����(�Q���y���q4�]��m�����[fn�!y����/"Va_�����RKQ�F�N�Xn��Lg�W��In}t0E��]Vx��J���+�f��.--6o���ЖƱn�cHC�ث��$1iX~��)�ͥ��l5&
wN�[Sts���j�!>fm#K"u����dd�I
�9n�EIl�2�e��qXJ��@�iV���y�&_"7�*�oh�+GH+KI�Ը�s�%)Bl�B4cC|K�����Rd+�F)2�7���
� 2�
З+H�'�|v�VN�y�q�*Ҳ����5 ��T1���H�d��׭^-.�J�ɜ�d5��>~
|a��y^N��H���[�#g3���@`�f>{�DS~q�j�K�C�j�uvEb��'�T#�Bv�c6��F�����2�^���;MZE~�I�O���_���,����3؊_��a
�Ѝ��j���TE����*�D]�&+���ׇ�n�����2�����%V�9�+��ԟ�l$9��*a$���YJ�u���â��Xb�����y�@P���CN�i]�B+=v���tq�Y2ZW4�k����x��d��E��v�:;�yX�%;�ao�wOj]8%�e�+YPgĚ���Й�J�^3�,�p$������E����$&�����cG �w�ᯩ�=u#� 7�tR���4c�jݶq�b����|5'�Ʉ̈�;�`[�������V����K̸1ޑ�H�1�]h��me���Ӵ>�ṋ�ރuđ���t��X/c���o^����u�V̉
f�o�y�Ǩ'�Dü��]H��tq%}��'c;�*�3�s��7�����OA)1T}�DcfU5�K����Q����՞�����b���N#�)z��˶qp�G�K�ē|/ o�$�m��vۻ�Ҽ��r̹��X�{�ғ���W��j��7�U��ڎ�"`��+��z���)�'ciK�;��
:[�2N6�N�=$#������X�zs� Q�EDP�U��Q�� �X]bӢ@?$�e4UA��U������+��q;����X��q�eL5��52x�Z%�J�H�B<�G�!���UI������&6�ٌ�!0�m���/1�ѝ�%�Mݴ}R�ݧx �aE�0Zt �0�����xFY�8J�q���{\xX��=k��+�*����Y��:�j�t�p@땀ϫ���=,h%��>��N���%��c��rm����$�jy�(�.��K�8nR�����Q��0w=����&���� �������>��ѿ��A��Y���U�E���_�	d ��,f{�e��g:�
4�(����
e��Z��-�|HP&f��t��q��ؚu��`�䦼���	�m?����O d�_�^ݎ�K�b�o���J�v�Y+�i�u�;���h[k�|Z��!������������1ӆ�Sc�,�;ʒಏ�)��͌'��v*i�O�zDB |�H=�Q�v�+`╊��"�cVE�e4�4�����~��ŋK��3~uj[T���2�bR7|+��|J![2P�V�Dt���ܵwi���,��c��pᣇ$;��qP��j�}2h)֤�k:)/��0���V���p|gE2M��,�:�:m5���i)e�)#	Am�ڣ|"c�1���"�?��DM~�DЊ�2����x	�����=3�?�U˸�ZE.7oD��;Ҕ��M&L�B�["����[�H\�^17^�9�0�V�ҰA"`�cF圽5��hR=ŏ��Di����� ˎ�7�'���[k�u;�F�Z���$(��n������Z���\¨OG���uw��]n���0���@p0�ǃg9(�yV�tɂ*Y'g���h,��t/�J��>L�� ��9_5)���p��-��|B���e��D��Ț{e~م�����j@6�k�K�3ᐻ�b��'a�����Z^r�=5�4J��frv�/P����z0݁T��}�����F�m�sc"������v�A�^͋Y�3�|��G�T�b��֓q^��"�)3�<b�G�m��Wq�
��o��\���J�YTq������U;oS�� ^#�,�;Ȯ��	$S����� &^�9�6b��l� 7��w�s�B.Zm1��;�U��T�	߈���(Y�sZV?���U�,)���ya=�P�h�Ӆ3��Fw��^½P ӑ�����%˧�[�ְ�ǝ����"j`��8�#t��m�L���D�&�v
�1�X��i�X���0O��M}?>τ�.+�ވ\X�+�����V9��/�=DT���������@aK�0n����'�|pÅV?�-J�`�FH\��l_I���;���J���V����S��V\('Km+1��N戣���iY�3�d`��bYZ�A��m�Uy)t���A�B.qE��#�H٨����@�a��t�p .��� �M`d4`b�� �hz��ڲ��ď�
�����D��p˘���	N&����d�#���Z�BOHv�N�;Sj#�JD��x9N�����y��Ё2|���o�W>:�P2D���q�Y�l�������1�U*]_(R@���=p"[P�R���R����EQ�.q���)��h4���h\T��[�W^t��C���G�D=e��ъ�����H���@HG��:w6�J{�HDX_R�W�$�G�i��E�1���$������5�B�A;}@J���jqg�P>�g�����9��vB�X+Nޙ~���Q�K���~����T��\l]�*���z���~�.
�Y�f�h=���d33�^�qHv��z�?��zb/�#����ќ�f��8O�(QA.�*���a*W�z5�i�2���BnP��������8�틷bBX5���ʽr� A��g���x'@���|���O����@g�� ϛ^�Hk��U0�_��5@�5�˩ǁ�y�b+�>�]�%�Z�}��n��y4��eϫE}���+8��90��lў���,,;H�=�-3p�^/�jo��Oe�Q�e�D�	�]$��]`5���*�}��%ԥ��)Vt�F$��4�Om �00�Z"�ʥ.c���I=�d��b�'�0>.��%Sn%�_���xܔ� ��`z��`�w}�!k�/�\�A�	��	/l1��5}��"�q����\�a�N��~�����"�Tda`F�t���-&�`^�y�UκG=��c'�|�A5��-A�c�N�D;F�����0j���u�"7֖9<Y����G�AoL�P�BXi��ۼ�jh�� A��k9Ԯ�����lt>n�,;}"�s�k��oʭ[��x���+�!�.!q[�^�|;9\>��Wq�ƪib�r��RcQ�ɝbP��NU���5��َ ;�4�CQ����#�Pv�-&�w�-zD4��U�����Lz��X��$�W��=k�z[�s����	������D�������ͣ���^��>1&�����}��nk�H�]�R,̳��"���Y	�e0Jk�,�tՈ �j�1�x��&�3&ւ�?E��x�zr��iQUR״k\���y�4 b�༉"z~�"���.�����O�H�X�`=�r*S�=������5�� ��Ù]���+:�M/*^T������*ߞ:��}q��y��~ŀ1&��nxtk����U�':8���0t�������C������"8�Y�,����;4+�Gsu�BPi�8{{臈s�/E���0�nq���ȁ��F^�<��ݪ?�_��i�"�u�3��"���z!�?�+(׀=b�2�;�ub�� ��],�>]�n�ObT?�&6tӬ�kR_ܒG��w�3�Uw(���k�TvH���Y�+���a��IH�6�,g��^��d�P�8�0��~�2KW���<;�D�}^�ǂ�::	A5�ӳP�l�/���=�g"��C?���:<LG6�w��=:i�':զ��	�!�r4t�V��,JF$9�]BS��������������P^��[U��ֈ��������dW��#2����{�ºR΁�<��s����&1�P���?�gk~����|�8i3-��ݟ��*|�F��AŚ2�U�$ɰl҄��!S&B�C�6Zq���ֻT�e�[y�N�+���C�-"�p���&p��;3�e��j��1�K�@W���`����������=�E)"�K�ꨅj|dE�N��O���=�V�r����eQGvޚ�)��0��D�a�%�{��x���@E�X���b�&����.�H%�SQ�.�̃��Q���si	H��X�?��i�Z��6( 	��YfY��UTQ�dh=���Ψ���^�v����d�����۹��S7�+px�3Lm��*`L�B������px{��I��D�Z��j�F��U#!]��j������j5�̄\-D$A0182�К�N�W5�V�,���dN���n��_���ڧ�Ozz7�ݺ䌾�Ѯ�N�v�o�+3�okm G�b�Z+S.�D4:��6RqEm�Z7.�ϗ�i����h�I'ݨϒ]$Q�D���|qw���M���|�S�IH/q�C���H��vvD6���vW�La,��#sz��HH�!�Es�.I?�N��,�
;�Wo��c���l���FGDt���i.4�9��'H�nw�L8�`����A!񚽠��|���5v?�^�+���oi�z�yBj�ayF 6N�!5c��"w�y 們Z�9o���4�xXo��Q�@2�Fc��VGPk �E��fX�h.;�$\��3�����Y*. ���"jV�oР�]�f���0!z�G��#yR)���+9�r��JM�C�E��O��w����v�~;�i3qeQ�~!��6� �g�K�����|��!J|����Uߞ��Н�>u���P�l�:�z�0�tٳ�,��S�)]ւ$�_���������Ͼ6�6����b���hd<�Um?+"C��IxH��76��d�|���J`�e�b�^� ��P������<��>������#xP���"�_[��ؾ����#�]+;6�Tx%���!��k�]^���}�C�����T�bk)#��Ͳ<鍩o���<�!�?ۼ��-IbJ�@�GH�+�C��a���`���\,搢;�p��d���&�s�؞.�֟�������ˆA?�&51��LIWº3�`=}3����e���o2��|���v����LO��N���Ց�xKR���f���Q	���C�����ډ{�C��T�e��xo��%�f��M��zu��rq&�ZZ#�I�yV�|>*e�TpxLĵ|f'j�w	�N��k�V8q�)<q�5�N���M�ԕ�A�4N}��[ۄʙ���)����f�E&�9&ƕE ն����+(��u�����dC���~�P��t�7+;dy�h��-�Y�L�s�7m2�ë00�4�4@�W����K�����TT}��m�F�r��f��7�Bg�/h�����u@�+��S�@������������g�/����F`r]9�* Q2��P����YJ9��~R7�_N][ Zt��d������.ݻ+�v�y����i� ��B�$��HTF�6�, i��aHv���
-6·O,M�T|��V��2��P%����.-V
��p� ;g��}g��wS����6��Q�0.]^��1��J��~�J��<��M��q�ڠ#�;��S¥��\�RB��ֿ�]l"��/���^��8�����\��k�C�	Kkg�#�R�=e��0�qǰ<Ð�.����[�g�bx�_v�6�W�F'򨝥�=���v|�gB�R/�5�?`���-�#5�4Je����pн�*�H͢�������{�N���P�Q�6]>�+��}}�����t*�)�,�5�9��o_�1�"�H�T��_R�A�놘�®��+�Ĉ�y�Bc�o{VS������#xd0n}����	�rn�kS>�aa����Ot��?9�t�������J<,��f�Q7�7�׀���Z�O�s}���ꄣu�w�
�B�	fJ���ߑ�f�(V��|��`�j6�W���nR����y���]�����"����)�`��$�͠��;�g�
������,3*uA��ƢFQ.�pW-J�9���QCD0$��9�Y���g�u]��c�]���jl� s������v �/2p��G\�XI��f5�A����|�%�}��o�L e��C��h�t�mz�E����%��V�hjJZ�W8ԏe�:��$��?�Υ\�e��G�Rs��3r�/�/�=��B�{�)g�ۑ�g �S�j�28#9�����ܭA�xM]�cw�sh�N.�^K~����o�����n
&�=N6z$���/H�>�^5m������\�����𾹡���榩�ϊ��n�P�:?��s8�u��|��!�,��{�K��X/�]�_ S���x�ڞ��,�����S�Ã9R쯙?�ί�NDrH���
��O#i��H��o��Dا��{��m����6O��԰@�����#��D�����yV	��GJПj�-��M�ZqO,Ҟ�ࡻn�_'
m�ſRE�h_Ra���0�b�:��pǄPs&hh��R�um����b:ح����5���3\K�~h#�����`>�P�|���7&#��n7>��| 8v�]G#&>׿I�S'.���������r��j��-͞����P�^�~f�.f�s��%9B-��־�ܭ*'�X��C�`��~˒26	Z0�o�H�/;3�f��Jy�y����4�7RG��ҰJ-ڳ|**Lx�8��g�>�~_A��W�q��Y�{l/?D�2Kx�x�K�����ZWa!Gn��#���M��K�z���Z䭖�2�K�8�ñ����BF~����.x�f��5*ogѶO��oq�z���c�$��G��P$�c��ר��2a���eSQFᢨ����[�2�E�m�@�����`fЍs&'qG��W��vz�.����m.O�(=�Kt�t6����+w��Dq��0'uZ����Zj+�����
yX�$�o�gA�l�l�Ԗa�֓�@������Nջ�QseO�x�ϒ��ڒ�5m��{�^Hy���`F�=�!4LS^��}<>���>m: ��Д�B�`�ǐ����\���ٝ�W��j���?�H�������7L1�ǣ����WA{n�c�rt�k@,�Hq�E�&���X0�Zi`9�^�RU�,;[���s�� �Ⱦ	��b<�M/Z���u(�[����s�IQ����Me��C陎��]��b\���]+Y���ޯ���A�ӛ�%)H/>m��x��eVV8�WiX��a�h���Hd۰u�_�w��P-�>�����;��5n"z�(a3�yÕ�I����z�"$M�s�M�:�A?O�AS�Xa�%Ͼ9,���+p:W\*��/��K���Nű��&�����~��(g4���&|z��;k�$������o��u���?���¬���"�����\c�z��i�`�׶(�5�E����T-}G���k	�����ɞ;ՀP�B�p��aF��v���5Mb:��'�<�S%U?��ODuG�YOCS����K�|&]��pM׶�(�}�2���q�6o��8�J��HB�0 �Ș��y8���09w����A�}�1��|���N���OT=�\ju�4(ق�	"pŸ���b�chiAro~��M� 	J���B���?3�b�d�ƅg���Y�wH7��+���F�@>�!��|,Ha����z&�7_�A��6�x�h��,L��赗�$�w4�� ۚ�ԉ@���`)��X���L�v�ێ�)^�^9<s%_3o�ڲ�n*��}of�k�;���#��ʜ~�rR+�I��tDp���^^�q��=t5<�ꦙf=V���]��S
k!<ǝ�u��d1�Rv��}	yu�Lsр�z9����s	A�
F�������� hI�82���r�p�����4���#M�hL�ӥ	�@�sU�J�PH��j�lIbYq��2ϰ�N:�+e��Q�s����v�Y�Ƿ N@ �=Z����)�JNTD"��&)�\�,��"z�T��ӹ�EF/�&!�C���J�o2�M�D/�,/��wy�$,U>��8Fm��m����sDg�ɸ��&�Mr����z�v��?]7yD�4eO��q��
	K�f�DY����CF�i{�һ�Rs۳cK�P&~<���<��O��C��G�Q13��XL��
jg�~�RS�/��9�y$h�ľO��	����-�Z؟�ض�,n��3���F,�i�]v��c~�q��oH��l�@�n�lV�\�h.�*������3�҄�z 
]J0ޜ@�2�Q��օ��v� Z�B�זmd�հz�+Oy*�p�:�c�� �7:,��91΁�$an�����@J�
��Қ�#N�lB���*XB�e�����k=Ǡ�� �e�0��w��s�)���P�oSF��R�5.ÝG�1��<�[����6Jc,@/��4&ճ��� MUE�!|��H�	�E�9&"}�O��,���|3�x�����.|1wV��^�����r���{u)�sA�,K��a�:l�+@$��Q�?���u5��k���"�{R�i��>�(�Ǌ��/"��+�8;�< �I�8�m����ʄ^�������UuQa6�K��EL�޶��-7�C�ٵ-����^���Dp��3��ÄLy�A����1��	'��\�-����hf$�	�\2�%;&�wmD�
�l"��tPz�#Y�\�tT�Ո�?���s����z/%�R�׬�����9&�o~���g��o��.�qvv0�8�C���#�3|�X	���xH"b���u�!�ƌ��_��Z�.� ��$�I�"K�G	]�7�ټ��!r����5�B�je��I�0F���)T����"�g3�1
(l� ?��!50H�X`uC-�������m���d1��̼ŉ/6�t�ʸ��J $����uL!��X���zݍ�=�����B�C��#�I���+h���j�v��
�5E[�?�)I���L�-� P�P�+o5oN���m�D�����1���͋};�y�+:����uel�G���lZ>Bj���Pk���iq����o���s�D=���^��FZ�A�ZxC��|o�.��b��r�~e4r�����S�%|�/	��?�|!�3�H|������+����pr~8|]+^�C�%ܬ~�$j�|j�R�('r�r��sC�Nb|�����a�7�E�+VAn�?z���1H��I��i=>y�cd���<�j)m{c_�d����#!�����Yr�����F'<W�s�뷞�����%�j�팴���S�y �J_T{�qiI���5����Y?Z[*�r6����Wԉp���|R�y����x*��������;Y@�_9���8)���l�{�-.�4��|�	oe�#1O�R������!P���������6���!��c}��>\R̨Q�;��/��|�����v
���u\��o%m{Z�j�h�
�2tfr��p�i/k*`s��(	�ED���V�W��{#!&t����3�zm�*_/�h���`��!q���3�å~q�v��ᓪQ��E����E����d/ �~�G>Zf>��;��_���b2	���@)��D�$�W�_�A�C�\/�N7}�nO4��u;B�fnh �h*ۺ8���Q�Ly�1��e?r)C2���$�Vϛ���=��.�f�>��q/1f,�ƛ?t?����<�����i�ArB�3Hф��i
r5r��@
},��]��l>Z�ƣE�k�ܗ�̼��.~�������q�pi����'��%2��9�ڂ��� b����O#�Q��ˆ��yl!��*��N��'�{Q�	V��
3O�Ntb�"&���L�ܜ��e#�JAȋ��Xd4!c��v)tT=>������Г���۷���T6S���>���BQc��	�M����� -�_��!~��dڂC��+Ӗ�`���兌<G�;�Z�1�����^�]�qɲ�Nn<�EPmox߼��0-���D<��w�����!��}
C
 �m�������uk.RY1�����=ʲנM�r��^�3�n�̀ �g��� ��aw��R&	i=tA	�q�����A���' 9D�3)J�߯'"'���_"�M�ᡴ0 ���-��A�\qK\��i���Eg�b��߄|�<�C�W�n����;)<\�s�����{�V�0"��XO�8���R���h����E?fEQ-Ij���7q!��<
٭g���ŸG��I�7D�=-�f.HR�u��Y��I�r��������& �p��w̶s��j�1����p��\Ǌ#y��$?2k���Wo�"]�r�`���;/|�$�4s#vz&1��NfD�@��S�42�?лZ����ڏ��=���k�U[���*��v�v�����N��&��sh[X�����'H��h*%!����k5�C6�J�P���[	t�`(�'-�H��g���w�̗,/F��5`f��<�!�Щ{�K�k&H��.�ͯ����X�@<<e�Q& W�c�A�%�)��	^S��M[�3(`�N���i��^-=�y���ߖ���dk�����g�����e_`�� �V��)���-��� �
=�)V���3�K��[��,#ګr��yh�����u�s�$����$R�?*ˣ`YBn�y�nхd��x	�FWL>t����,B�D�iI�G���� J|H���:�^��g���L �a��ރ�'�a��bc�)v� C|1v�z-����9t`�`���.5�+�:*�N�È�te��:Uε�O��5�$��Uh:X��tT���P_��u�9�d��k��w�P��VDr=�Dc��'�ZԂ~��B$勘�k�-������`n�X�@E0~P(�Y��H�?J|��?�qMn�����sCZfK@-/L]�=��8����=|'{m�o쟵H[����XS���b���LՖj�K9HoC'/T��x4U��ZX1�)u��CI8��O,��ә����� �:�
���Y���tU��ˬ�7)�q����vڈ�e��Y�{�F�/�!�Sﾴ�R2E�\+-FK�˅��rj�<Ū���R����sC���Z�I�Wn����(��n8�uzlwA�H>U ���-�Qj#�Am�������0ڧ͊�e!��ٺpI��h�pTI�,3%���,����?�{��5N�ő7/��8%a�ӆf��#�½Bg��?�Dv����h��#j��A�ɣ;��#�!�XMv����9��\������$u��a�==G�e�И����Ƀ���0K�g�Z��#_��6�y�m$�۬_X�z�F�L��ѫ�O�-j��0 Mc�������, ���ӄ����X���1�e�F��dHHw��7��4k�oTҌ�� 譊�ޮ���P�s;�.�w2D߹�h���(O���5�F��<u�� vFaPrŭwX��m�V�U�Ww�X Ǚ��+��S~S��y��:�PW���T�X����إ��,�U�0��;߯�t����\"�#(px] N����b��1)�^�u��)-`%�^�֢��!���AD|������usD`￧�帎<딵y�F�`��յ�q\6�����?>��H�I��&�u���C� ���Ŵ<ܵ���#s\7�=�l	��e�=	�Ki��*���}�i�1U�ZV$҃�و�*�c��|��Z�5�>MZQb���-�l��	�Z;�S�,�9�ڞ������:#[�q˄Ƨ0`-5�"Us� /���VI/�.�7i�,�OG�6/����6׽T$;�ASO�є��%`��
��ߵ=����u�wS t��T�!Ö���`X錾zDL���"3���z ��Q.��ɓ�'P[�-���6Q�T=Ӝ��s}�Ԛ�AS�'ZP3��ZP1&8��m
"���Y��Gz�^ִq��E�l6���eq�������_S�'&�� �WF�P�՘�����J��:�k�Y@�7�k
|\�}�N�({�ܮ�bX��k�n[�Q�f�����v�+ ����"p�I��M\9��y����J�1�Q�Q`�Ai����0�$s����F���k�5G%�U��g����:�)��/�b}e���s%g��5��\8t�mC� �X*GvY˻�s��i��]�ZIg��G\��A]V^�s���� ���~�a���sE� ���?i�~���`Zd��j�]�XQ�u:�o�7
�UW�w���c=b��,���#f� ��d&�Q.Q�01`~w���k�����J�[�Q�sUxE_yz�w���R"A��v�I|��|�}������e'x*��~d�Rտ�m4{��Z���Pe��h뻮m�g�̒��9�S��5~��"�9��SE���>�!�ƐQ@4�H}ŏy��jY&��+�*����6�;�F[M��zZ�%�������jx�N��Zo�"
%W�������� ܺݵ`e�S�er��]�籣��F���j�ɡX���~:`��5�s���G�4d���	������!"t�������%�Tя�_Z[��+�8O�l�-�^��2�_;��낡k��H���S�nY�A&�xd�H�#��&� ���&c5��[���q����`n��S�j9P��K�j<�mQ�������P�����YR����c��SY�[�2q�h鱷�Yѳ��ѨO2��
�%#�ݪEk��|�U��<��ƀ�;��_@ˁ��� �2����?O�z��Mħv��tt�y,���N���X$ ��p�����H��k�����AZ��l�˒���"��q�\0�TQ�����o~�Fm��\I�t��t��(m`�7��|5.�x��b�3��mN7�%f�TE|y=<���d묇���3^c����	[^��Q�O@Z�
9 �V���./�"��� �R�W���h��]&���do���{þJu�ߤ�~�U{�����7p��7�� D�4��P�14�B�ɦ3�[���;ĄKV�+��q�EF����5�ȯ�zp5�8F�{��R�?5��*��=\�SU���ʗ�����bzɩb�u���^f��_2!�-w�`!���^Nu���Y7�����2p�R$��Ϊ>=�x�=p߉(`Ƒ��~�M9�..��+�a��_!b�������	�YK8��e�B�}�����P���n�#��w@�Pt�b��$և@ߵt�ĉd��E�JJ��4��m�0i�Sݕ�m��bM�i� �c'x@L>�2p�B�T�6�m�&Hs2�M�a���#7���S+����Z������\*��#.��,[	{�&n	y���{k�_㗦�	[��:���U�Ck���(4i�G����`f��Jw�Ү��|����U�77��������]!a��d��ڏ�=BŨ��pl�CDd��A����S��M˵Τ6�EІ���_���ͅ1Y���� Ȩ���?�q�?�=,�V�q����*B>����G�̩�͔�R�vu��	���]|��g&g�w�[H(;�۶��(��p�����)������m� �)��E�2G�х8<S��ظ��]�	����i흓e� �n�b��5��r���#�>��K�.l	��^㼋���-dJR�S9��Z��~�w��w-�a_R�� �ʞus~*�=h}~�? `�gB,d;��:�h��off�;��})�[%�.Ƙt����v�A��w�d
&�=��8��?��E�'Z���h��"�o�Z��	��`��Ni�E
Ƣ&��8���~�E���*䄘J���Mq>��&>�Ĳ�V�2����FWEk��vz�9�vIX��R��#��N�Xˣ��%R@9�9��,[���@�v-�i�i��5���J͠"o� U�����kI �dH!a �s�M�i��_p�K��"-)_��p�dB�H��0�愇��
}�%Ba���� �F�����ԏN՛]�r��a�ҿ�ކ-$��@�4��4�Y�>��`q�L�I*+��{�b�#7}���$��Vm��X>Es7ٹ�zjc�;�m��;��z��(�qľ� �X<JRL{�ߞ�Dr��
7��I�����&E��
ZZc;��b@*�j�$p�k0+7����A����b�}�Ś< ���)�<d�d��;���8���<��+�ľ_�Hݳ�]oܳc���R&��*�6D�t�U@s@��m�}�W##M�i�:��KB���_�j��Y����;]�W��^^�c �n�az�P:����v�Z=��FIn4�\�q{��������y���*K%���3Jӭ�N<0ȋs���J��ctG��D�	�Y�Q�Ob��b=0�QI���~�8���ߢ���	�!b܌�5J8�5���SM�[��K14V}#n�&49<wu����rt�:C�		�)�	������9 ��l၄��Z�{��y�����9����Pn�U^m�د��O��[3 ��e,���~Yri�n�����4�6ɣ�R�9��QL�L�Um���ߧ��oĭ�-��g����f�8#)�P����xk�tZ��FG�ex��-�v�T_0B@u����WРghh�T�seMF3�e[Ow�y_q<��Iu��Zm�����07� ���%�q j�ݶ�7�^c���*6��y9g��M�<߯�.�F�40G2�F4^�4Y��~�p����2ȶ�,f����%*����s��h�H@���	 ���+�@�4Ȋ��g��F,����|�,��?e̙3�	Olg�9R�Y,o��*����@��q����u��i�ĳ�z6T� 
T$­>�z����[�D$�y�zB/<>��WVd�<�&Fj�g��f����7Y�Ś2�t� �e,}Eo�Nbe�h��k��fQlͺ��'ܩ��,���"�F�#�Y �=E �E�c�dp��5��t���%&����0��sAC�r���2	��
�N*W�׆L��ҷ]�j9��cd	�}�+sā*�<�NZ���+�e7��#�L�D��H5�������>��~N²�=Җ��:�w�%&�	�[�Q���3f�$�fA�N�ϕ�dz+O�����Z:_�;*T� [ү7�:T0&R��
��@L�u�x��hZ�@�p�ިWƵ�$�?j���y�˄���L��B��� ά �,����Ze����c��}���
s��(��綇O��70+�xݠ�u�M��*w<�m�jꩺBK� 䅭D��Y����ʽ<8�Ef�U���6�$�颜��<��dD��D�g(q@<�'e�zp�Wl�	q����x!�;���ڳu� L_�9N���@��+|�8m�����}	9=�BA0�yۘ�7�o�g�Q1�q���@���(�I���;&QB�� &;��w�a�� ?,Ǽ�W�B��W�`��cg����;pA���V|Y���}�邬�;��SÕy�B��a��:�i��RЀC�n�W��MAo��nDh� +�n�I1�>�������ܿ��7!�y2��qwa�2*��a�{SL�����_�'eof�9)rm����X����oW�����|��U��5q��>��KZ+ zJ����]k���ȃ`�p����H]d�p�L�.H>�`7zF����dNB$�&� u�>�L"�s�/Z��}_��^V�������%K�Ѣ�_�]���`Ξ��(�e,FD���0�G�giq�ߑ���uLJo�*�{�<�r?㤏���җN�E�'�~־�� ���������y����	*A~����gԠZmq@_�X�)I�d��b���E�^	�o��.?i�>����V�IOe�5�@s�Ց
oFf�e�0o��)1�z�l8*$�KF�&������!^�,��[��O;�U�ޢ��S�~P�0!@���pl���Ѝ�(5_߈.l5=��xeH�ŏ���ylyl-���^p��썙�LVP�y
��xz_'P-��AB���y�k��S����:.�P��YD��J][9d�%A��'T\l��K[���O�4)����i�i�u�+ڨ��z_Ѫn����r�*�eiS-����ݎ�L��ֽ�z*�*�z�n�X
m�)�X��>�|���P9���'�#M�e\���@�sf��.Au�,�	p8�bX��C�쓷0�~x��q`;�?�/
� ]���Vf^s��V`Ia�QWL 5���fm~"m�)��l;�� �v,\�8&0��>4����i߯�4-}�
�R�w5��s%6ꃬ�x,�r^�
�� Hq_�O覐�%�]�[6eUR�o��-L곏F�a�2�&�6�(y$����
r�7�f`9�Hy�V7N~�b������K��x
��4zB�m�i�9Hq�o�FlY�����h�R}8֖�c�5\����\��)䊋��R.��,�����R���19a	�Ge�y�Y\�C�6�,��#>fS����l,k=�)����lV1=����a��<��ĶVS����4�O� W�eeoP$�1��_�K����Ӻ�!��P�! �YE�N�I�	���h?�coRi� �$zD�n �W������],�,�L%v��$����3w���y1i]�E�U +�SUB2�ݬ�$5��\Uf��3/3#~R��)�4E��Q���\<�|��� �$~�`GQ$�V�,�@z���E
��̵�8��Ize�l��YL;d�)e�m@�ZZ��}��Ҭ#[�:^�n!Qdh�pZ͊3����Mł)�	��j����A��ƍL���5�q�����.���1��ť��g%��뵒�#�����},�f�����m���ߗ�v�H��*%e1�0��K!��ޔwT���v��`a�i�B.�)��LYb0��718� ޡ�!�� |t?~��2G���
o^�#_�����C���#n1T
K�V�&/��M抵"$R��u�ٸ�[A�f`�TP;��b���eFu�@�uŧ����<��V�Z���[��Y��*a���n� "(�N�#կf3
BŐ�(I�p`�DA��.������!���}��˃� �/L��]�&;�в��!d��B�)�P{�o��[50����%�����z�cN��5hr�Ă��U��i��bZ�<���֦�jD����=Y$ے�5QmÆ�rѽ5�9*#�Ǽ���K��h����m���;BHp	f��Z��3�#������h�ϲ�O�CfN����>���"����z�?��q���bK�z0�oXUO*�Nrg�#O$**:���S�d�A�&�|M�	�ڶI+�!Σ���Qb����ح���[��6v"��&T�G���(���%�f՗�_�	G�ƣ���Q����X*�S[uX���Sð��H�cj���(o��	���[3*� )ǩF-(���K���'�xng}�kH�}Wʫ�h�4hC1v��/�'�Fw��^q&4B+�xd@0���Q��ڶ{��m����b�ۆ�GS^e
���Rx��}�.�3DQE�"�z˳�A��C6�+�� [ƴ|�R��B�\��E�x�*Dy�Ͷnn��Q�6��b�Fd��߳5��H������%��6mRŊ�^� Kh�O+�}�!�N�V�����<J���Zh�������Ϸ����?K�e�OR��x�t}��$�U���g�R�Kݫ�U</.��^�,���)?��k��f1�^#���u�N¬��)+#����p;k$>()�^��˻��ZK�1٠L���oX��v�̇�f��F�=v�'�[?iD!i�/���X�!�X��[�镶+���?p�B�q}n����*-L7�q[�I��6�o[x���&P����L�Ͷ!z��et�m��mdy�=e��Y�;[���_���U��܉*�%�Hy83�@�ٍ*�b��h��M�6Y{��+:)�o���-�`��֥ *z�g�C�����2��!{߇,���
��Ǝ@��(���p�z�X�%���	J!���� �A�����J]��V-�8����$K��8B[�~b�f�b�ɋ����nV��a�Jz⯭Gzf	����6���X����r��4�ѕ��&U���A��A��xs-lذh�������~��Fvb��:��E�k�I]���վ\.�Y�Q������-�6�:��3pD�h����� pKZ�	^|5c
�;�eN�d�&�\�|zn~�ѵ{'����r��?/��!�x���(���h�Q͠z�E05V��\�.��J�<m�kf�s�4�<����Znm.t�$� �0�d��;;(�ᓁJ� �.����f�A���,���M�ї_���V�$NH��#�p!<�\����_�f���ij�"�v����e��:*i��;�d�Qo�٘��w�i�}ڡ�gd�~�EwvN\�t��JE�вpJɶ&qdi���nKp�!�m����-�����>�w�(H�m����/�����-f��vp��E8M9�Jwe?4�Q��м�r�kp���G�~ ��X��4���e���
������ŷ;	�,�<EE'�R:�O a���g��C��5�tZ���z���iYL����)�k�l���Ї#��+�룟���UY�+�A��n�s�~�����\q8kߦ��w�9G���$Zq<߾5�QU[�i��.{F�����C������5���A�K&8��,Q	��.O,��N�hD��^Ұ�p\m6�<+��N�=f$�.�e��x�qs�z.\�s�n�	(�����?F��,���zh�+H�as|�'p�3�Ǩ��"D7�g��
t�r���[�]��(%?�����^CoLd=7�J�ϑ,�y���QޘNڿtȉ'�Z4�5����~3Y��\$+��2V�a|$֖����Mq�)z㿚Q��������I�lJ$n�WC^U��U�]@c@w�(�������Z4��0�Z ׈��,%�0���5��<���v 5���b�^)Ҝ�W�e���Q�4L8d��E)F��Nh�<�<w�j��%�\QO)vwWHi��a;�>�[�	��7	�uq����6��D�����)&�*r�<�ZĮ���/b9�����&+�T�E��TG����چ�R�[�<�Jǀ$�o�Y���8N���D���{�{�|<�Қaq|�<P�%��+�'�tjq8`x�XV[�HuM�z�Yݤ9/AF�����)��hP�7���P1)��C�_4��M�w Tu�fr�v��'���-����`��r��.[�� '�N�����(u�~��yޛ�E1% q͗�u�s��yv��Y3�e� �Nu�A-(�m?�C-.՟Oxf���G�S�Hq��~a�`�`z��Wۨ\���[�Z��(?<�y~��>Ã̑9��*���5�k�<Ġ�apk��\�'˸P�y/!eD/]º�⹿��U�F���5t�Q�9ǔ�oh��Y�k���j��&�?W�!H�](��n�F����ʧӧ�S.C�92c��X"�L�;l	����<���� �&�����.�9���bK�06���!E����G*g_�S�L�]$������>�`�k��Wt�eF���.ml����۟�:��Y�A��^���WVh�q"`؍�;�]���M4M;��'$@�=�S)�뻦6B�D�q���L���`z���bK{J�p�^���1~�6��񔚊�ޮN��Ct-LgB<b�~N��X�k�{�/�����F]�������+��x ���)�ˎ����ѣA:��SӸ�{]3�-�-�����)�y�;�'%z��s&x!�r��iI x�[��ڷy��!�0O����AA�B��"�3�H �U��	�<)��G�Ď�����m������'{��C�H�7�B��f�����6N<�|�>+�^j��v'7�5�-,���� �Sc"1O=Y�hݰ@DD��>LY�}�Z��+�s��[8K��!�W',�>أ��D�݌@hM�M��� ��kz;�8�C���?@�%�V�sr��/2 �%�\nU}���D�96/'\�;,�F�D���ɪ��V��sq��[�b`���R�H'�u�{�༹a�n����OΖI\��P�����}�����AK�0�[%�����ٱk(iF�b�hzJA��Q˪�p�cL�C��4�7,�q��Q�q[�l���U,
�L�g��u�1���?�=���=�Tb,�x8|���1�j!��	"ӳs٢�N%�㋅��n��f	�0��=���b�'6�^6�A�cvIJ�~�v,�}�!8�y덙��q�Nv+�=ʕY�7���v��|e����'����b	{���\i�$�^�{O�5���\60zT|��Cod��7��W�M�ΰd����uԜn���l\(J9�o)�.Il��c	Ւ���v�&Eq�s9�����	�q힡T��۫XӀb ��G��|Z��Kz(o� ���V#��'̅� �1U�K/ԗ0�����_�zT�L��xςX����w�3FX���];m21
cB��QQ)[lZ=�0lH_Љͮ�๊%�c�����J�����6�[i�h?ρ�A5���k�&���D�O��
��y{�B:�XbG���a�d������K�]�|SH�Z5tf>;k$�*&�",m���k�G�
!��	E��@`��&��e�V(/=��S�\iLN�-MGRjf�L���_��տX{���)@���ӍCo*����J!�����o�~�5e��^4�N�qc5*$��W*<3����չ��mj3�
�Ě��#ܥ���xh.h��g4Gm0 �T�$畤/ݵ�d��!���^�$�ϻ)sU���p �M��Rl����?�OM/�?�G�1�q[&)۽�����ށ�o��=�\5VsN��Ÿ��~M��6-��t_Lt�:S��(����<�m�FЬf�ue'�胐a�;����M�8[Ra�ꥉ�)o/C�(DQ��$D*���͟\���),�o�>c̮�#���ܻ����"�3}Ӵ��b��������Goz��&;L�����y
��Y8(h�O$g�*s%�f��W�(�z5*�ݱ��Vwg��E7��UH���\[ԍ{�H�|qiZ)b�3�7?��-�q�3�$b�d�C� �<��(���wP@��ؘ����N�N,ڨ0{����ZVçC.%�䈒�Z��rW|�I�0w�|O�g�/'�*�iq�}�1�`m��f83�g'e��̖�=:U���I׉w[:R��*�k�M=|�	\G�F������0�1}�Ц�J�Gb�x)fX�V	pk;\/_�4�%�'j�ʢQ"�Y�)�`;�mQ
����@̽p�.� r�a]�M���8�Ȩ{��+��&뺉X��"aS̮�P�?0~�3�&2�J�)Iy� �lZ���/X����#C���i]�?�Rt[^�D��5����9���-��� ���r�N���)��ƨ�F�"����QTι5�ӟ3�p��:P�o���6�ښ�$��&r���yaA�Y�M�ѭ&��y9�Ά�ǰ�)	t774=���h/��\��_p�P���s��\�I�^�h�PS*� ��O��P4�������9?�̆�EQjN� ���r!5y�M1�]���4���i�n{��M��P�bY�\JV?
�5�[������h�]Y]gAS���f?���9�r�J�=���
.X��J�K��;JG������6��!]�o%x�.�	QM��VAy�qTT2ȣ����L�H����t��i J�Qg��m�6�}I"^�o'�F�Q	�Y�Xw��Q���%|��d�U�*�*>��<�Y1�5��{q���i*8���U_9�����V#�9HSVdIE_�7ಆ�u�
�4��衧��$���nI1�
���ؽ|W;�o�9�Y$���V�B���8�F�.i�� ��y���ury�̛�9���^8	�ʾ. ��ƚ5*�;��/�����Ze��&cm��¯̱
��5 #=�F��Mm}��ԍڠj���Z�b�י�v[J���0��K�C��	0�!l���xzC17�O���F���&���L�sQw�h�ph>��d���>� ����������OhS�����c��W��\�I�7C
�<`�'%�%-Pܗ���	*��'tºM�L�Lۘ�.Xr̑�є���f���{YEŽ��Á��Z����^@�'EqV	����I�\�t��B�8���������f�z	a���gf`�IOY|C��=8rHsUҦ(x2�y-���}'V�ר�Q^o��Q�A�[voA���j��#�a��=��ڊ�Ӯ��x��!�3���\���7�"�tC�RM�3Я�t�SIwiЊc�3еܬ��%��g���^���jW{��n/^�����дnc�a�5���~���.�o9�ؗZڎ�H����`0K�m�Q�{��f�K���(���;�\�7^�/��!;�� �
�w{�ߕ��˸�0�P������ߙ%-4���]Tp���^O���b�ܟ���h0���f��V�P2x�J��l�����}��� �5B_�>�X�{�"���<�u�}=UC��x�E`��+��/&W�+�1��*k�	�Z�U�P�l�4g�f���^|�Q?4�)�90(���+A����T��a����ږ8q�B���u_t�P#ɫ�b� LFm6�vI��9΢]v��_�&��y�n[+F�i�l��3i��N�P�d�P�E1}�I�tN̘�J�@����`��@�\J�x��*�/�zb,�u���ࠍ�-r��T�|�!i^wb��3���R[�e��� �x�Y�����`ˍ���<	uE�a�U7���dP�t0��|/���ø�Wo�OOi~!�{��)	 ���w4�ͦ�t�MV��[&Z�yTj���mH<.�r����	�>O�oْ�P����)\��uԪ�$p��ON�9ʃ٥ib�N�5"~�A��G:F����z�m0�i�&ň��==���yh;�.��q7��L��&�e��q�����ݼ�j0�TU�{�_'�A���ďT'Є��oj���6�^�,Quw��I�+��+CK��m��3Q��[���?�����Y���/f"\������?���iAմ>0N��iJ�bZ��	��LS�.��*G!v�zW�P�15������]�=�<~#��r5r�Ç��\���Db�d@�2��
=K ���f*X�b4>o��:�����l�h qA#|+������t|Pܤ�Q�������yw���B�ǲ.��٣:*���O=��!(�L�-�3��6�Z#'�Po�/[]r%��z��Q�P5J3�O�Z�Ŝnhp��Gȅ,շ;,�p���c�4}��sI�5g1\9�����ϴµ���G��)�'338�?�����n�RJ�#�W{p�`�Dp<���1�&��׾C>k3"�O����Ͳ�;���;|!���b�\�l�ԷFe��d���bx�W��L�7�+1�q���v�Ȉ�;�p�7#�g]��̀��cĻ���@X���,_������B�nh���=��gC��d�������<��*Y�KN�g�/�M	�F��,��T�p�y�a�ɩ��u�������F�l��Ҝ}-3<A:��xZg�yܿx�0,�������ӣ�p][��B:�|/����c�*������)�/^s�K�,�>�F�C��R��p��${h�%���Mv�F@�5w���u(K4�]?����0;����K�M�$��>$Hm������]	`�*'X󋯗%o.�:."�Ns�<r���*С�GF���d�	��ch^�s=��|lb����k�,��w�dk�D͆�|�����5D���o���`��8�Lo��05[ý��״�}�����p��"ߕ��a`�-�BX9�'\�T9�8��lD_4�a���av*�8T*����S�kP��7r�'xT�\u;�5 �g�Ƒ�Kq�`F%��/�wu��1�FJn�2�#T����m=�0�m�'i������;�U6O_'ǧ�4��V=ta y����Rra�'�G�*�%�d����z�&`��7䯟�� hCv }�h%^7_)�>�b�ܩ�-ild(~�$������Fo�n"O�\,�����t�ng[i�w���Cx�����M	&4w.yJA��v@X���n\'�cz�Y���\aFQ͟S;y����$X���
x��۰�FYd��b�ٓ�-!yk����ӓ2 ��7�p�(\fJ�	�%PB��L�H۽"Y�ظ�����"��fF3�ǖ(�
ː'�2X�,�S-�N�4$x��]m��fXZ^�t
7�AicVǝqx̟��N^��)���su}�U��Aؠ���-C� ʓ����M�<����}('6G�W�q�-ʉ�6�-?��,�A>���B\�8�>(�����<<Ț�X����M'x��;g��Zt\��1<�|�^���{�
X����Y&Ó��c�� ���
K�8�'���w���.G��Xb�3q����h��E,ˀ.W�� NK���N���b�Մ��ߦ��L����F�C�[f}>��੩J�v֖2Zpa>�]i�D�A&��l��g����|gJշ��s��tY@`#p+��	ӯA�+������k�5�:*gh$�W��&ӂ�&���ۗݥ	2F�����HU'��{�ٚ��Ya s�v��$�B������$�UI�_[��%N�7[�9XqGf�*<�
C�U�3��OX�Ō���Gr�eUJ%�<6vC܍��4��a�£��8�J��-�3�2p é�Z:�������m�gnT�I�p����8ҙw�4��7_.��q��dN�?x������;��kjP9��1��"��n럒8]�"Y���G~�#U�[�I�������KX���Tn.���)��f.�G�O���f*P�W��v�ίUO>��Z�#\v��i�0�}�a��(�����[j$���ͷ֍�/�`���h(t�}�S�$3^7A���an�xP�8Ѝm�^�00`S�����Q�ا��M����VD���_dF�\�)֋n�ຳ+�l���b����vrh3Uµ����ο#��A�օa`G�V�b{�p_�i�WCo��=.��歅�ˌX˛�dC�1qt��Ӎ"V
i�b���٬�N��z{���QW�x�"���&G=6�́�M�wcU]��K�kh8F&Bk�7�,P�X�+9��c��	�kt���6��nGE�+=!����Ļ�^�0��7ҶQ���Y�]���D�j�1z��y]���CI@F\J�Uaj�@a��H F/ס�z��CV����ك�֚mb~��Y�w)��i���p�����P��̺u*#c�х�\h�wf��;��ͫ�V#���M�j��p�H�?���	�IVb?D������V���QI��(�?��=�8��Zqd;�G-I� ��%���Q��H^���"�?�����
{%�$,�h��� d��Q��#UѶ���ڣ74��"\�{x|����qB1'�<�=����L�QX�m9�1���8{|W����)t�)���R\����Q�f��c8=%dB8 ��8
.���ƾ�4_؟��v7��D-����zXs~Y�gڕF�/���a��>�G�����.�Z�`��=�Я��1W�0�����)1����;�qCI�Iu"��~G4 <���:���(O����ye�:-�c����r� ����P�U��1�@J�>t,��$s�W���r�[N��-%GQ�T��c(��B��}0��H�۫���[� �~�ԇԐQœ��5�\
���+(23!PF-�C_�S��Iճ֋W���kux�W?����K����Ѩ��4�¨S�/}���4Dյe�V�θU�v�
s�>֨g��(��da��LA�G��)���b�R:(�K�b�����`Ѣ�5uD*	:"�Q67����>��-�U�#ن6����4$FHj�g����h���mFR��i��?�ˎ�'���>��V�@� ���3j"z�W�<^xjKi�����3��u,W����Pk���9����{�8�����5���� ��`:ꍐ�r�� ��\+H"��G~���"*�[}z���`P�n���v�	�!��q�Cc��1�ޑ˺��r�݋o�KX��c{�*�%�tU���˺���D�f'i�T"��TY��o�O��7��d؜�Fړ��E�Q�Y�o��� ]��2���s�]��۔ rTϦ�����M��:+���O@�BF@������tp�
=b�g�Ѻv̑����}��h)Qk��Ž�x*��&�!-l���@(��8c��/�J�3�)�`x���E!����y����Y"5��o�-���o?OLy{a��fG(:����WX-�BX�V�z=lqg����c��j��\�l%x�k�mLD�"�K��_�(å�i��Yh�+��!k�4�C�.20 �ʕk�2�J,�nu�S,��<��ɕF�(�lw$����p��%�1�P�جxBP�t�����X�ة�.�|6�Q���0N�ZJ�ɶuֽZn��Y(�CX��ɤ�q~j�(J��H���3n;�ֿ����H�������xY{IiC0����m��]�����w'�Hړ�����Yڳ̖���+���Ӳ�lbY.����K���Ф�X+Fj �Tv&�G!@�(�~�z�kk\Nb�x�06������T�*�Ȑv�1yX���쳁$�S�pE9���~2��2����T�٭	xC Ub���9~���L��
K�TfdZ�B����~���.x�"��tr�H�3@'�ku)�\���V.���2Y�@���*�[翈T�����U���l����W��>��y�]\��}��Z3n�f:�ړ�;s'��Ċ��e�<n���u�x�U�sȡk�d��
�_�4X�����f�?����X�e��8\Z��p@�J���/���xĬA#|	�A��mQIf H�@"�7�����co%�y�0r·��B�������6=�������?.����cXo/�V�]`@/E�ScF9_T~`D8�U�"��8�f�l��?d�L%q/�i�����9B�N��-�N�����a��& t��'�D�p.��&ш�Ytgn��`uo�[ٻ8����ʈ]$���/�1vc�����u!�L�ʖ��ݗ5�ہ�����w�����Iûr.G�uO��O|����]\XG	�م���h~`E�6Q;
�V�zAlV0j9�zɌ߆ނ�gS��BP6�������U�w^�ck�V	!ܝ;����Q�{O�},�kB��9\��hK�_�,=�JU�ηEe&`�v?np�#�u=��{��^�G+�ǋn���T5hXj;��ԍ�3ڙ��[E�:�7�a��e����B�x��竉-l�υ#���o�dT)��'k"���~�����{>�_h�S��xY Àr[�3ѕK*���gT��?�AK���J�Sg�I�����?�R�6s�82$i�
�O��g=�B���s-|��!��u�7�� ��-�<��$ ��y���k�<|��JE�2d�������%�)mR�e�$\�EE�m�ܕ���|du6�Wj���t���l���h����&�4�������� J��B�i;H�r��yLI�7;�����~d��0�X��f�b*zi*M������ '�E�*�x;�M՛��@1K��B��o��D��-�w�\/��z'J��(�w��~/-Z��փ9H��B��d�R�������%UL�R���ͅ���5h}��1Hct �T���ҭ�.����i��R�(
=)�T�Q-��zPwsey'��W׶l��L�K1L����1?��`��cQ|�v��p�P�;���_c�T�3�fi:��%�:RM�R�������S��v(.�ht�`w�g�l��ǳF����nˤ{S1� g����ɶ,����&�Y��z��=�%���
��b���+î����-uK�Y6�9ص�������t��1�'����"VBT z��������BaK�V���R�j����E�^ۘ'�Bs.xw�O�v�b9U�_:�m���_dv�P�
�m��܌�b��WQJM.Ecڴ���^����#��O5i�3��b����s}�"��{�>|I����<�(����=�ꐘ�OU�ӅU��+��]%u?��7)���X����$l��bWK���� ���Ws����t��6���K 3y�� RX&.?� ��l��~��y�y����3p��9����G?pS�V�L֤'�(\�|��89����g���`�1O�������	�xz�\���"� �����ɡ-�w΄��ů��ae���<���0��[�����@A�5���]��ա�I8
xCi��Uu�d�� �x�!��.ǌJ�6�Cєu�R�(�	F�s�S�1AnB>%m�5�k&��䅠���y���� ����~I!����.�rJ�u�(�Y� '�&�|lU8��I����D��ʡ^�l�o��GL�M�����V�u"SO ���ک;$;r�><�5���&��)���)4`��:��6ޏӚb���j�����</���{�uS3m'���5O��Q��	��^L��u�u����\�uz� 	�A��pПf��
���0F����ĒѶ�_͜�/��ύ���w�@.�jAv�������
�T	9�a-�Y���+V-h}�3^93t%x7K#��1���MՄ�G��:��-6�S#V����FY?�R;Qɡ6����%̔�?�Z8���ψ�о2b�eV�:7�`#x���7��a�rF]
�G^��>��]������3�"�g�4 ��U�w!�����p�:��h��%���@5%��J:��[�$��㔓C��E\�^ķ�:^$9��s��,3Uƺ���,b#����rL"껾(l� ���Ql:FȾ��Ns~!����(g�n�&f��y'�)�I!�~�(v�C��1�iX)=��0�N��8Y���J�AA�x�\�o��y(�����	)]9�iyuڻ�gq醑Y���	�^�([cjv�
TTO�rcz��4��'>(o`4Xe���j���aċD�3C�2�*�UiSSp��<�3(d��9�[��D���M5�y_=n�A�,��v�Q|�0�鱩Y}�:���2�n��.e����t�
Xcq�dF��me� l"�-4��l��v�L�B�>C��p��et>�p�n�����T��3���Z�4�e����&''>�D7�U4^۞n�ߝ�H㵻$�*�0-��6
��Y��ЎT��~�o��)��~uC_v�7dϨ	t����-S�������9J=��`X��kE.j�<W޵�,�x�:e��w� ��q�gгbb:1��K#�.E��=��U�WGs�K�\�O�H����C��1[�G�Pc1[5�9�m;�IvH��=�6Fج����4Z�x���0���I�C�4�ͱ�J����L󺦕������m='�����쑕w�+�u��千��T�&[f���.�tC���/d�eS���B4��p&6e�I��t�{�3�ҠԋX��ɂk+䢀���6�j�m�7��xܒ|"y�5�6u+�[y]�q.���4�ʹ+�v^������|��>C:��K�A$3���	/�wz���S:~;R�y�����u?0.V4昴f�nY��;�X�6�d46n��68�D�UF�����24Y��3(��H�#��D��&���<٭*�t�Jq
�q�k�/�֨��Q7�@�&>6���rueL��#blB�ϡ��TŷP�}oU�b��6�jZ���<j>�;��%=;hV�ᬐeL�Yyj�4�3��d�4�����6�������s�ˀ�wo���[�����'�W���Ǥ�v����9:s:���Cc�'���Ob���; 'pZ\�h�yCf$���s�ճ~]�H�;Hr�%�[
*��d�π��8'��j�_^�m�?�P�? 눲m��?Y|/�$˃~�V7q(�/q��h�y�d#�"�8�f=G�k��Ն;R�d6��� ����c_�Gk�ňZ�7�f�>�~�$lLY���D�"M'[\)/�ɨ�X�7�֪*�bY��e�@�N��B;���d2�/"o��7v�o�/��[�?��W���n�~�G�V���58 �������*�N�J45_A��zC�ւ a�x�Y ��s=�E��,|�yC{9
}КY�t��Y�p.PL�䤿6�͗kR�<�@�g�;<)��z��pJ(�һ0�*��Vǝ�	O���%�Z,� ;��^�����[|4z�:W(� JX��D�i
�z���
&�Y��ߖ��BHr���F���;G��6���my>c¥���K���@�Ru��hl95��~�1mYR�����O,p_��bBf6�:���8��IS2��DX����-��\P��f���Vjj�R� �|��L!S�&�̮C{�S��t|�{�	����Sz�ɸ[��_�~����������a���(e ;�M��Y�mObY�]�02�����XO�qMr��YP���	M�yX}䟾�6(QE������~|S��n�n���¼�RCo�5���S�\�d3O�a�*�iU�(?f���^I���7��l[���8��{o��ܢ��Րy�+�W���S{�V�:v��2�~�3�)h����j!G�R�"J�v�;4��T�ċת�%.+�E��@<�x�80�T:��埠;;�����^���p�[X��"��.ܰ�AfśK�"�P���<@��>����r2+�]���%�R�[�*��<&�4������T>s�3���1����h�?H���󯟐Z�� ���1�bN����U�}�B�ޑ��(Q��C��X�iZ_�,$�����zA�������^y�j���uM5�T��Z��.S�}�$'B˅��yW�gR�BT=G���S���MX�x�yX���(�X�_RUɸ�w�#�*����AdM{i�����X̏�L�cE>�1�2H>��� (pA�Mn^���s�)E����$-�Jp(J!���o�Q73K5��òT±�$9D� ��hVm(\v&:w�	^z��B��-��Լ��+B1��)����7w���5��1�~��DdVnע_)�!`&�����'���%�Tƒ�PLb�+��E��f����8�xdLn���-��?W��������Mr(^E%��q�*�Ş�\��A�@K-H�����b�ǨT+I4�,	"��[���fS�E6�_��S��*+M�c���@HK�!�κ���������c��g���X��Fd�A�z��"�GP���1q�6v���gp�j����)���g����c�+]��=|R*�g�ُY������'��W�P&���0�%���A9(�>9�����%��mY3�؟̈́l�V�4-�!�� nh�Z��#u�pH��6�L�E�:a�0}q��`�^ 3����+�N+����3�����o�"\�Q��WY�+��Q�<à�KV&[���|W�QP��� �{���t�$"�0�V�{	Y��&����l}��>>�,�bcq	�U柲���a�;������~Ay�Uͭ�!�L(�5]S�	���m`�p��nEy8Q���n���_�qM:g�����VA�����&}ر� W1�-�ƃ!��S���w�~��t2�~N���)�r�#�'��W$�S;���������b�����4�Ġ�4�Y0��U��U��TؕYk�RM*���~�=?�aOS�?M>
Pѩ���� y��c�2�=̜;�2�}��zM[��KA�IȘ ��UW�B������.;׹IW�3���zD
���Rh��\w�e���b��e	�n$5b��tV���zհetes@r�r�Yi>Z������e��%�b�����s���9����aW�:�T l\��Q�x�£E
����w5��.52�z��������p�h���α��QB��O�ZX<;h�n	"��VN?9����kv�kG�-�)�No�i(E���f�p��Уn�n�ل&��������sG\tzb�Z)y$�-�F�o���5fU���-��r��#���� C��W3��,��H���͈��Z�#q�<`˶tTY�F�.W�U�卼Է�Ёr��Uo��GXhҨ��5���QN��7k���J����ZR9�?u.�X����I�vا|k���ce���!��Aj����,t��o���,�4�,�FgT�~T�G�Z��S�^#��/M���p����J�ov�	)DǢCR�eP�D���(�:����UO�P$��׮޴���z
��-Zy�Ie���j�q��ܝ��� pb��8u] Fj���- �0��u�'�Jb+.3�Ȕ�9%'��i<�C����QD+���x�l_ס_�&��U���՗^s�:�|�l�U�nJq��V���Y���׬���b�Bx3!`#_\��ósudK�h���+	�=?}?!������ � v��:���]%��8�����ic�Jm���K�����'�qg!�lR�t%��pHN�q�-v@���3tM�,	fbһ�Q�/A�8,ᙜ�[� ?�̡�H	ރ�$�o�E�zs`<���l�O��b�����c"@��`�"�����$L�ݲ�_�b�Z3�&D'9✅T?�"�e���s�N�g��a)�H���l���<��(i+I�k	A��i�Om\\�Q����[�ʠ�P>���	���*�.}Y^��E��d��^5҄U���K� x[>��hh��M~)y�ײ��B]����Ψ$�L���b�Ȭ�z��w��e�,�L[�Ƈr��F��8 O`DO?�7�O�vT5k#BY�x�U!i1���њ����ҠH䏯�sݍM�&�����A�_��x7�@hAѡ����_�����I\�s��#����7�e��2d��䰀Z�jS)Ҩ/�]�f=KcI>V�<<�"M�
� ;��Cee��H	H4=N��Xn���Փ߫"�_]N�J�Y�=��i�[���;"�i������!��//�N�:NZ9����:bT�PCj�����W:>>�k�����N\m��)$�C�Y���ua���ސ)�}�Q��8�>�������c2لw!~y�a���y|�2�g�s�P���<5˵���6s�0Z*���v�n�AAƭ��F躒��{���|�le&�[��׳f�<3���)�����PXͩ Z�F��N���1;7U��)Ig���������@JE��9�{��F(��pӊ7	��<	�p�t�z�9��0|�ZAA��nᶖ���C�Wv�.�K��gL�x'(�1{G*�5���y�)ш������1��ѻ\������ SqK���4\551�t@ϭ��r��	 ��.�\���,�h� Y?�wy�4��﹈���t�*�U��kC��FU����6�$.�� ޠ��0&T�/���tUt~�/r/E+.j��tZ��pC�'N��h�'s ۃ�G��8�C���V��2��DW�ϥ�{.3zo�ל�9��5�()�m����#Lۢ�~x�d���ӎRLCdU�*|�����L|������br�B�q}lQl��"�L��H΢��u�M":��&22�&�mR�S�|�3�ي���1JGW`c��]Q�5m/�B��K�#��.��W�J���S�V�a�c���39&���Aͣ��: ��B�EVQ{Q�� �#�E�� '��S>�>��d���1:�h�YP��Gnc�!ĸ�qT���-}�<���f��5���?�r��#K�K��w5hW%�S)��ҥ2��@Q&;	��T�sa�̟��-8
�|���k�¥�r�8y3�p���]����eeCQu���rf*�S���t���x���J���13z��6]��f�"-R;�<@�<���>%�,��v��}�y��C�ж�.��}�K����t%̎M��7�0�.����_�7{D�$��Ǩ�g��4Lh�w��)!�39m1+��Uk��)�3E���)�	;g�jc���R�t�P��{�鋪�7��H�b��?��Tf�� ul~��@�O�A��bߠtRQIYc�@�7+i{R��#��V'�H�wH�^��5��`(��_z��p�L�̣7OP��J$L��(e�2u�;�Fhtd��_��"�]z� d�@���s)����@.'ǉ?�H����έ���	�U�l]�gm(����D�����Gб��z>Q��L���=@םk��xZ�ݨ(17
Mu�m^�ز�!A��TMf����$��	(1`�P\[�q���4'HT�[KÛ�Z4���c@a��\��7c˶�c�\�k�E�i��<B�3��V�?���3�I�EB&7!ɡ�]����]P��Pvj�<�E��� nmRpה˕��F�vؖ�TfT��M@e����`�t�〻r�S��`����T
iW��6����@�t �!d*s�oH{�\s �aFX���p|$P�Z8�_hӒ���Q�|!T�8W��y
v�*�j�iO�䩶J��f5Y�ȣ���\t;N�.W��*�d0�k��z���/�§ؐ�[>� UG<�l%��F7���9�f.)<�{"�1��Uʶ�R>M�V���X�Fn;��ˎ8���/����м&ȻF���=�j�$��S�]����?����.Ob�P]���wA)/A�~ՙ�xӜ� d �I2�|d����K��:ƫ��
M�n�5�i
��X���SΦG��#�>v�"6���Y�������<L믂�eѨ���1��P�|q���4���y�~
��_k�z	`�ftގ��G���� @�U�A�=�r�3҂���-1����>��	:��+���ݜ䐃��,x�A��?dP�,b��<%�� �%�;�0�|��.�E��8�-�ǢIB�����38�`��w��\`eq��ļ�x�S�_�̱�B��u����Zf��
	���K��-|t��h}X�T_r��3mAR
���S�Ȉ��x�r�S&E F�	g0".L2����	�{|C�_c���ۜ��6D�KC%h������u���������h�i狼����8�ti��ɴ��f:@���b�����WuA����ԣ-w��3�|�A1���Fs��]�y�D|�m���-n	��!a*�S73�Nі�(��T�p^�<=������RЈ�R"GL3i�;��r,�n,�,<>O����#��x�����`�՞�EI�]�î��'N�S��BNlw�������C��g�/�N�ͻ�7���Nm�֏ׂo5_�F"�����z�X g��}4L0��AX�=F�%d:f_!L�M~�蓸~pϡ^m�"~7ΐ�j�,)6$�[S)��1�Ijua�IҬ��ϡ6�*%Bs��N�P�����θ� ���A�Tu���N�6'Q3쾿���p��3K�|hC�^_�,�؄ݰ�g��B�1�2x�f��n��j`S&�y�Fe���7�7n�F՗Ҵ~��XFFd�C�L�	65�z�1-��ɟpBW��(n"Hd!}�(7V���u�Z�g,,шAz�A�U�w��+]fi�Ի4l���V�ؒ��6C[��!�V���_f�����[]��"*;�&��P��Y1�Ϥ���K3��z𚾜k)C��V��1M%ts�Z�9�A~m�A��������2���}����j������+54��n)�vH	�#��fMbљ�C�;m'���P,�Fa���*,9@��q<~��ö���Qf+�±	�/R%xD�E~�n3K������P�`4��Ae���b��7�K��D��CӋ����(�xV�����вۼb-� JA5��F<��M��ZD}6�_��x��r�XS�����0��؞gR�8����p��M+�itG^��̞���&4�P�ӷ,]�{r�ë�� �R\�����m�l�v5
�
ɡ���r���� ��3��m�
��D=/���w���aC���[Z*��ר,g��NS�
�!�3*�
��8�Vװ��K���U�� *����)�X^ه#����QY ,�@�M� �'7�`���M�S~��F%���@���c����3 ��d�3�@�TגD-�&w�i����T�sX.�͙��ýf` ����#� �+�D��*�эB��]�-�B�P�b�Hk�^����l���]!�9o��o�Y�!���y�w$�� �;#�ACB��& �#ҙ5w�`X�XMr8�k�$����r�!�S,o�0��B��wߙ�x��e�:{_ED�<`ƾt�����`r_�	�JKv/;p�:�
�y�S_���[S����@cu�\��I�W3ѯ([���N3���~���H#��V�����k����Ġ��$��j�C��X�A����;� �=3���^ �P�R՘D���[K�tr�7a�Ï[��N�(��7�u���*�$j���/
�Z�WT����:�7&�U�ZX�u�_`mz�o�b`ƣ1������mM�=G�^��2e@^s��x-ʄ[Q�Z��4K���Bun�G���\��)v�r���4/C^��!����ײ�T�項�f����Xx���c퀗A$ �pC4�IRi��Z�;(�6D��m�X�5�c/��մ�����ڳ���M��l{�K	�Zd�G�lm�����y���GQ�Ӊ~V _����W2��!h�իe�(���Wfw�.�o?Cg����42E����q0>�}��|�L�bM� �R�`�?$��u�;�X�U�ƙ�2%�[�u��C@�4���ܹ���wi<�tE��Oט���T�$�����
�1eʕ��V�`�g["��21qs�~��M�p������b��!/�g��u�ʋ@6�F��O�^��~R������ц#?�CTUs����PV�Z�p����O}�l.�1G(���쮧��ER	�*�t�{�`�LdZ�fVI*�)��&Dղ/�*7F�Z���Ĝhh�7$�k��B�f���S�бҕ��A�ZiT7}b6T��=��c��3MMD콑�%�p�A1�����<[l-(cz�3V�ݱۘ� s��p�g�-?�`��+= ۚx����e,ř���r�1륔�lMиE	�Kئ�bW,.`ux>m�  �-�w^��uX��5��ghu�����J&0"��J�@���n�"�f؛<#i��N'q�[�׿;��(M 71P�c�
��h��<i�l.��#	�)��b�z�B��ut�US�[?%��<��ӑ���J^���e��;d~Cl4Y��v���#���^&/�āܗ��`yY���*�,Rzڭ��ϫk�q��L���Rw�$�ɋ|��P��?}Y�(P��Vu�b�(��1����9P�؇w~:����sv+���Kz�	$&<5'{U�����hm4�MŎ(6�&j	��6|w����0�Ƞzf��.�����Z�,,�D2��!H��N!��݂ŜNqW��C�5} �����&L-R�nM96p����W32����M��qQN�Z~I.��`%25�rV�ʝ��V�e���ߊ�V���~﯄��ܼ�R:�	�<z�'H�O&�t\�Q��{?�<w�"p#Z7��Z��,n�"@�H��_�C��F5���T�1"2|J]�s81�W�պqT�����j�>��q����*�*/5q�w��y�zJ�������Fr�T��/�YA�9Y��	�i+,6�.�@C����{+|��ZKT*��OТ��w�Kb-� �4ˬ[��]�z|i�W(r�M,�f�m�T�
���*;���8+S��q������4V��ZP���k6����+ ��"=�'3������� 9~Qg�2��J���h��HA���Y��O,Lļv��"��`�N���(�-K�<�w5�m�/.�W��u�/Dt�l�q�/F�j�3͝�Ib�u-b��)<g��:�<�S�-�����dh��ក�iL�E�	8��������b\>W�m���e��4m��6L���t[oR:��n}��:t�xMw|4��u��;>]�)�p ���������:cVH��J�����)�c��\AFX�eQ�,ǉ��J@ܧ��*��?O�ܡp�nk�����T�Q_�����Xu,�I�E�w�n���}�U��D$���2���W-�W��{};�5~Y��~?��^Q^Z�% �Y��Eި����7���-TH��@-��,�������L#�m_�)���k�䣥GG�r@�晀�2-|#6��GC����,�U
��d�{m�v}6:��3/;�1R��NME¥�c�ǭ�2-����f�<x�Q�����'���f+�r���h�Vi<ݍ>�x)���CUx��{&�_�q,��,}˒��s��d�ƭ�zÈ�(�C�_s��]�"RS�׬E���S�uwh{����\3����7����%6�r�����a}6R+����MK!��x���WS��2�&�?jk�[��wڠ5�e�~�Մ~5uz�Wm!��q��X�B��w��P���e�K�j&�����F�u��ځ��5��\N����
w3��)T��Z��
X&؋����[ju����<1L�fZ d0�ݽe��k��pצ�O��~3�"�1~E��Zr2��U'X|�cR�+px��(kɥ��f<�kZ���C�;�ǋ������Q�okȬ�l���Q!��A�W��J�6�G���B��1"N�`��s�HJ�-L�<���L�g�>�8J��eypapX6���F6��<��Q����8�ߏ��������k���fyǠ6�nT0���{��p��:6�(������ǂ(��#�����Gh��~k}U&�O6C%z�VB]G�2��sO@og��yP�LE���$c�e�{?(*1A|?T�&��~�Xn\�d��[c5�N՘#����jk���+W��LQ>Z�P�Ԩ ŹM���l�)��=�\݂��!��s�t�����{7-)m*5�k�\����4��)�-јR��2�M��bZ�,\SJJ�2��}�W'��00t�&9*x3�����&�R1}��u�4G��Mx�q���\Rηs�����+<���RA0ReJcيhk�Z��:��n�,(�L��.�?S��HHw�}�R�]���~�k=tg��W��ܲk��x�[�[��k�Q�}����*[�n�'�f[���
GqG�DP |Ի����0�Ȕ���v���*���\Y�@D�u��K����ؔ'�hR�,̗'��V������ T�Y�z���[�Gu��)R;�p�/��z�B1,��f�k����A��bA9d�'TY~{Iz��I������M6��|�l$�;�?п�Z���! ��Ŵ/Ūf�)N����l�9l�I�8�#a��_�s���2i�����W<��9~���&l/�5$d���s�4��)�jDV}m:x���x��77#Pq�z}+�g�x$�e�֢<*`�����W�i���H`��M^}������sÅ&�������f� ��s��L)�5�HTrH������ƚ.�������.����7\�θsAð�+KA�aE�f�����
�x��kr�%��$#��c����R[5�v��hrw�x�f���-K��H��u����>�[��WR����v,,jBvg�����(y O,�a)1_�`ˉ��\l {�WhѢ|��ub ;tk��z�?Bw�I��,����;�Ps8�x��ކ�p�꺣�����a����<�:�ۜ2������B#�9��q�9_�_-1� �[���U�9�ðE����ͭ^-,4�=E�����|������k���!,عϢ9V�^�5Y8����C����) XN�Ub6 �27[X;�͇������lb-�������VIrmҦ��ѓž��� ��r_�Cx�6�K���	#�n�����8&�&����։��J��YѺ��?�j��_��$��Sd������C��a6Kz����S���}]mʉ2*I��3�����ϊ���[�.ݦ@�<*C+��0�@���VdY���̱0���n�!�2#�X�lX��6�2���6�#y��TXS�F�5�|Y��;O��Fa��ŶSu�e[��9  < ��f�"�\y���Tׁ�U�!fƇc�t Nm(l�<�
�;]���{d����ot�C2�%�^��-Z����me�u��e�E��tX���>/]�P��0��YY�q��S�(5�%��k���ϴ��ǂ��	�z�` N���9� ��,�g����g8�n����I����c�����ٌ�cHmZ�W��žε�{(����6L4�˪HG�����N%ܲ� ��� �����%ajD�mMcv�%�W(c��,�xrO:CP��	��gu�����3Z��G�[8M�Cla3;�}�m�뭂�Q�7������ RRKyŒ�.�^�Rs*�]�����K6��.�"��$�!͂��2n'QG�8}"+Ѷ�f��[�ϛ�o0G�T쁛E��a#��%`3`T�FG�7�sV�е�o"-�X��U��k`� }i�o1lܩ���L7�v�n.^:�Õ���I��鋤h��k)[��æ�=����a�ݒ4����#�k��r:Wt]Z����R�<�'�;�]EN��pwj��9���7�Z��n5�/B���`���:�����F>�(��� "�~X#�*�2��o��a;�0������|Hh̪���A7�����L&�y|+���_1
�0�
��&{�,�on>fs���:/ם����7�P}t�`0r� ��K�8v8��,I�D�*�!�xqH����t!=#�Ҵ~ߗ/G���x�~�ɹ���E,��-k���~�2q�UR���{�Շ�Ao��;�ܡ��Q�����J*�[��ДC]O3pG�i[i���o�Z��q�xM�l�[WO�Z5n��i.ղ9�=�O`嘢xUϰ"�M�����M�$<��5H���޳y�	(L�����A˛�h�����/?ٽ}��_w�VA�g��K�$��	΂�"B?�
�ڎ�ʝ_JS�y�f�w3Mq��4�]�%vt���%������l��6���E{���UZ��{%W]�+����(F%tE��w�֬p��{DD���-���D<a��#�܇���f���K�D����8��Zw������>> w`����#I"�
1�iH�B�K
��d{�nq,�{��?se�e0��ɩ���D�<lĔݩ�`��M��ȶ�a�t���E	�(�9?���% �ь��%�!�۶�f����������jQ/��)�/�eE� �l��g�u;�Y�O�M�ue�4���������F��A�|�l�Hp`A���:�T*�ߧ[���T0{��OТ5��C<�,v>�8�m6m�8�w����P"��B%���c4(�F��t�+$�'��:kW6�����m�*.�X/�ڞ��;(=B	��R�xX������sꂔs�x-�Z�{7�«�x7�ju;��Q��P�A�}N���N�u��#�~x����F|
.C���[߫�ri6�i�K��e���}�����/~�s����:qi��&��'�DN�Y`)[y�S�a>�r�=<Or�j�q:2�d'j,�Lz��#̺����r�3fU��"ϗi@�vO�ÿe��]���5�1yd�,v����*>1�4?���k�u+���>�������T����G��,���/S{[�n�� 3!�*\
��D	�ɵ�F4`)����}[#Q�ǹ�1���;�(8V:ҭ���b��f�6(�jIC�,g�;���Iiv�h&�g-�K��X6�ѵ{:�!�U��ڶ�"��D[�F��i�Y��\1�Q�ޗ���)>�UO�z����B�|i�����L7�'���=�?R]�A�$zxV�*����2�y���L�d@���ժ�	�����Je��e�!����?��G����[D�,�{�M��Q�1�i�E1��x����M�����v���tn�+6mE	*P��i�99κ.[�����QO3�7gU{� �|s��*F�Ek��Q
�+��V0.�v��?��)8S�����\�A��H#�jWsk��C����"�Br������NV9e�s���K?{�S�m�����#�N�p���X` �ҍ��L�F)��M�Ӈ\�$GM�ʧG���I�1�ʷ����ݳ�ה �x��L
�b���+�9L�����<�Ц^[����c|�z������sE�`xF �v�)�EG7o�x̭������_��]+PV_0Q�����v޲Z��/�{��&�d�����e�E��4n�:�7ysU��i͈Q����m���~QP�xz���j��%+p�[�q�î�����V^'�h�[�A�1Z���5�
���_YJ�'B�<[�e���h�
m@��{4�fF�#ϫ�x�-��t.R�3]5x��?Nt*�."<|>����������ݵ��ݢy�ݲ�<D����ύ|M,%���!	{�:���>�f�2��,�ۂ_{�0��r3c�ɨD��=��<��=ƽX�3��L���?����Gq�V�\�!*ﵑƈ�Tj(K!�w�=��sD������5'I����%co��-�Yh�vT����y�{���jh(�[�[�|�?�/�]�)&�{�xP�;.s�d�-L����`�)���1��l�Ȃy���$�i�ô0F8�1�hKm��j�� â�c�B]e�ү�}�)�K�������/���҈�����J�Us�� G]8U����*|�k�UN�t�sY>T/�b�F������R����Ž�	=�A(����73�_BM<<��yE�>z8C`#ΨW(�d����(��n�����qK�39J���n�(�Y2�������l����=�$3<���F�2Sn��>�@[�b֧�L7��7s��Y4��"�x������e	�E��G&��J>�@�WN��n���h.'�b��m&�w��dh�q��Y�>d �~�%\lVL[�卯Cn�f<��H76 �x!Y�{p[�����@Sˉ�b�8E�5c��ʐ+{�s�_2�%�E �#�2z[���D���k��@ܧq�n����1�|�i1R]����W�{"L�Om{O��B>ꏳ�Ǡ��đ��n���e(�KSsa�J���	� �/� �j�ERk�,آι��ٿ�6�7ʂ+a.�!�c	.�I��2*?�$Ӓ����li�����֠���w��7���8x�s#�<a���3��s�a!�K�NB�Й��0�2��Dy�[��1F�0T������Om��墇i�
M_��]5v�<�'Y-g8>P?�;��$����ӤS�����FlGC�_��^�<��EIl���r�Ɋ�f\�[������0ǓkOq�]���Yq%(L�;�`�*%��i����,~}~���8O�#�A��;��cc�?%#�? �0�B��|�&� ��3y���7�(
Ż'j���f&ʆi WH�K��SG&Z����#U��	#$�f2��|ެ�Z��K���;����y}��")��qk��,�ү`"V�QGm_3Cx�1�!K)��>QT�7�'�օ�ڔ��k�O�����'��f�u�xک���tUICy���e��xD�KaL�|j�+l-~\�eb�e�)��֒�ԌOx�H��+����ޘ�/��Dg?J�_�/~a��� ��3:�,��lT�m�� ���^Oƻ���>J� ��6��LN���L?��>t ,$o�n&�=�F�y˲>M7 ���;��s��e��'��/uͳ$C<�B7'H4��֫1����mJ���*2\��u�R$?��}�p�|�L Ͽ�`�+�I�D�l���W�5������߾�}Q�ό%�N3��X@��5K8�����������������<��*�D���_*ʚN>���]��o-<
������J�[Bu?q?�©��:a>e4��ܢ�Ӌ��,�OxZI�v�GS0��_J<C�`��~� ��|�N�-��7����Q��� z�qn���R�����qI�}����{h,��@`��b��v��&y��6	F��![W�����5 ت~H>.ts�Hi����_����R���?�A3,�����`,�f�7d��/����d�Mv���;����1��Av����-��%�� �gNsaƎ�ьv�g/�)V����y	���.=��̋<��m-��7�hۀ��U9L.xz,�8�K1�O���Hmq���I�\pN��}mYy�i��h�ɱ�Y=A�"5nSa!r���C�O�X��Ҕ��К>b����W�$T��3s���4+6"@Kp*L4�&D�g�U�ݦ$��`";���E����zȃX���*�->n�K'�A.!���m��~�姤��~7X8������c5���p�+�b�'�e���*���K��@��[2$�d�NV��-��q��A��yi�P��}�2���B��I��j$��� ���"�Ȱ�.�0��TP�=X2�h0L6h���W�~Ŭ���o��	A�e�1���Q�"����?�3$�-�$i�{S֓��d������{�|]am�����$0��
3͜�����}� �(�J�M�&Ɏ�-ߋ(����S��h6eEF�8����wQ�����a�3�r87�C�k�J��T��Mh�1������4������*��Тk:]��Vf��FJ�D���7]k�5�APZL(=��uW���w@�^�͗���_��r�S�OaZ�"n��#�C�Y|t�Sc\�0 ��,�-.DOJ˻ :�񃇸�P'f�����ԗ�a� �@r)�Zh�q?�� }ECG�7��"V�&�g��:*!�ׅ�z+=��Kc!���9������j�G^�N�C.�!o'c�x�h�D%�3���ᢻ�)O��-��po�����s��+��*l-0��[�b=bޗZ�4*\ �DT���K�-�R,���+�"����9^�]�?1��Z��|nMx\�O�gjuK����}�&+��KP`=l>f��=,��]+C�l��F�����2�3U�;(p^lӀ���=�L�(��qͮ^!��Rg��&R�	#��#�ߺ7;�p�!1�	�ɾ]s��UK��R��@�@Β�NR���FQ5Ш�Ԅ�F9F#0����:�{&�R����I�1�}f<��e.\��I�lN��o�U�I�΃z�p&)�K tS҇��N!9���޳,J?�h���x�NL^7<��;�ŔU��ŋ,�TR�n��$Ph����3Z���NW1֡?���S:��j'�;i����j&3"jQ�F�I��� �5UD��'�"���� �N�2��5#�����؛B�8������&`��7E�����������?g�e�:-���_o̰_I��G�}2?I+�����\��;؆���^J3ْ���Np��cQ�/�E�4sfе9�����t5%_�'qak$���A�l0����6��
H=d�Y10�GX�dL��@�}n\�:�g�z���,?�'�tu	�u�U�r9k� �O[]�,��$f)�v�mǠ纃V���/��v@�e�
��~��QQ�����^Y�&��򔆚��(��w�2�L�dM�GCk;���(QU
/��Z�����$����A0��RVH�B
���'Q	I���.��2콚��p �b������;/�"�&�h��ʨ���8�(��AO8c`��ݐ����%O��'�1���.�Z���!�Hr�<���2�E�o�J��<>č�f��5�զ[)����2�`T�7n�,g���Һ9z�aIx�*V,v�TlkJɝ�s.@˘He�˕�����]�P�Ƶ�!ëqɏ9Z�������B�s���],������֊Aާڇr�W8�$������������ީ���s���s!sW-��U��=ROY�@�v�4�\Z�G۸�p~�7'��9$O�J�8���ΞW]wx�I�@��3'�f� ��ӵ���/)��G%0�+���V>����ɯ��ɰ� R�"�]��&	���۫O	��W"_�2��x��o>���c�khC��(<�Q�>/��U��{k���y����GQl�G\ȣ��+�]2[&��x��y^���R�>}���;f7���a㉵�TU�Bvs!E��Sb�"�ǲ'���Ѵ}uB�\n]�' ��%�w��4���Y���������k0�&���}�m �̋�q��lzR��VD~M�dY�TN���ۻ��i�<�ڋ����1�>��Eܕ����"x��ph�מI�"�Q���r����|�С�q��^Q����G֞�D@�被|H2�4����6��[�$8<�}fx�������pFi�J�)�Mrm1I6����`[��㍌�K45�9��P� c�G�	�ӻ��&[�9���NXi��^'��C��U$�<�g�����ˋ���DZ���j7l%%�H��n�ģ� 86��Bf��]��b+fVAM��/��,�ۑ{�����93O��&� �'���
F��`9]�Dt�Z ����<�q1C������_�"$AI!i)��Z��!d�+=s� lK6�ѷ��:��Z����{�OE�^g���r�+bC�f���&������Ⱥ�{��kС���d�|j�X/��R�����:���%���`	�oPtȓk�����E����ٝ���J,�\�Dx:��C�����vl}����2��=��ǌ��-E���z	N *����(s�`'Ϗx�b�uf7�Ab��f�IU.���%���)�ǓF���^ׂI�C|��8��/����/���{-K�~,��k^M�3���ٍ�\�djj?"�G'��o���eh�D�D�>����-j�S��u�s� �uR]��U0~<����~z�GQ�c+���KÜ�����O!'�U8�؆���Xs&�H����'olB�V�*(�z�uc�V�\L�AD�ӹ3��gC<}lp�4;ӵ����k��+��3��X�v}�4�<�&�]1����^x����Y�n&�"$����i�	]Nj�`}s�M�bD��c�`�y�����}.�#���Q�O����O��F��vW��F��m�.gZɾƬ�V�6X?�s��1Eio]��b�f�N�ڷ#%qȈ�����!SY/9��F?Eɤ�I����T��)l�B�F�G�E<p>F�(�N�ڵ��R���;�N�%�[W|,�����D_�>����d1�f�����}�\��w���;'��L�!���P�疺��f�_|$��Z�U�u>f�Z��D[g��hF�L�i8b�It,6(wB8�����z�/X�nw�a&��q��'/T��P�(���S���;إ��\��-���y�Nm���qG�	[6F�,�-��Y���[�Yϳ��R��~Ϭ���޴Kܵ��_��2���ǜ�>�uo��5�0\�CU��.4�Oɝ3!Vl���4s׷y��׭�0`mpb=���۽��D�X�i�����-��]J-�}.R�����ky�S���$�;�)��,�7��ǲa����Ţ���^ٸw8��P����E[���a5�	 WVGC�������vآBE5c���a�w/�c@��`]o;��9�����]�v�+�Z1�
���kg9�ε0{&��n [�
J�X����(7����Zhd�߻�W�m����ӳ���{��Fc� �Cʭ���8��鰥���C۶�"��>����;I�0�D���dE���C�3I�B���k2�',�Ԭ�p��H��ؖ�(�`[���Vmd ��toA�#��[���YO`I�#R}���������9��Ԝ�[ޤ���Ge����d�IL�s/�:���ae���k<������Ƿ!^�4w�} ���Ġj��1�}pD1�=�1L"�[]$ >
Y��wT�� c��<ϋ���)�ƨ�>��$�'�k;�G����0!��X�֧y�6�����OL�Np�v�**s����?�ٿ��s����e����T�8y�.R�vh�j�.W# ��)I|�OL�N��ʸ���ǋ�����/� �D�E����R���_fvAOjq��������e�ɿl��e��T6�D�}�0�\����_�%��z�|���UXV���`�b1�PZ���cܐ����c؜�Z3������#�>}̶7&z��S����b�ף��a��v���+=�^U�8�`#^R\�u�s��n�g�4f�n��r�)�Ł�4k[F�kW�q��U�kY�5�!��PEG�)�3п��9{����8s�P�ҿ��v�N �nD���*����{��\�y-n��(P�;��PFr g�'>^��:X#��Lf�i)o�j�+�É�=J���WP-��e�S�>s�KJ8��)W�T�ި*l���#`�?-����5�{e���$����K�(ʚ�@�6<�;,�,w"7O�� ����A[�Ad].^W\�=Y����He��-��W(3|ϫ��PǺ'RŁ���.&@]���ef�����{�:�Y�&J��� �i3\�ksQB����#VH�GC�CR^���ܷ�#t����r.�4ze|��L+�[VWA��kDP\�g��*���8m�)W�L�d�cIb&��C��O��eIo���3кsR���2F�G_���m�u��L��tt�ա���T����l	��G�R��u?q�86>p��~}�|�W����aLݶ�!���M
��Ki�F�N���;\ġa7NͶo�.����d�=�(�E��I�ܵ������AlW�����8�Xu��Pi%007�Eh�H�Ĭ孫߱y�31̪��rY�3��|�e�Pg��,��Mw э�yFY'P���G��5"�3��Ҹ�H�)ꌋ������Tz$�r�_�5'�E��l��=O^�H!|��<�p��f��P=��oU�2�$����N��70Α���n�h|��'$��]O\4
U�֡-}2~��0�<F�2��� ��y=�,qX���Ȳ�����}ڥ-{��o�AݰX��u�
�"�D�%����t�������4��a��r�Tz�l�.R�5J�=g�u����VT���L�9n�������q������p�\�|��گfrH�� ���"�͙=��G�z :춢*$�XT�%	k(O"��+�W���y6^`΁�<NH�Ɍ	�CvF!H�^bs�p(��L0Ѽ���,ξ'�2~w�Əh3������A����`$���p����3;8vǁ�x>�"|$i�ɠq'sG��M4A�/�)|�jsU�ı�����i`9��B�t��0ȡ�X�m��8�ԣ��8��$�)��Y4-�.��`@��r-銪�e�N�K2;n��s�ɢ�Jw�'�֡��"�7��mJk��h�=q{���T�.�O�zg:h$�V� AVU>U�ğg�y,�q�(���Ͳ��wL�+(x؈j�zMA�W�)��ۄDV��� ��S�:�L�~s:��zU9�x�8%�s3&!�K��ORUꔖ���q�x�exm�y��OΉ����8Nx��Օ�Գ~�8�S{����7dU��ЊIS�('K%��O��>��\�pq��$/��h��V�%�Y�Il8v 1I�/��Qt�C?��]���ܶ���n�އ����gZ�k��Ҏ�aÀ�X?��.�����ϔ���8��+������}q`� �g3Y�:*�'�y��U����"��5�S֥��{i���9e��3R����B��*X�d�e�@�K�v؉BE=��m!��v�6ܼ���,�*�z����K�G���T�,(�Ǽk��
ە�l���L���S�ƻ؍��z 	4����ſnR����'2{ݕ���e�����1=��+I�W�+��Ƒ�4����c��Ԅ�C�t#Y���W��������l��.@���QR_��W��v��%fht��)|7�&�}ZG�����G���J�YHb���<�J9nm��XF3	µ�DȋÎ������l@a�N��\�YOE�}�@C�@�o$�����m͛�b�p�bZ�-0i��HT��O"a�NhkE���������ĺsGJ��z@>����/�H��n'�`%���_Y�m��<���9I#PS��*X��N�r8��d��t S$��U�:�p��o7�&>fY-��i��z)�ʨ�XE��(�>[E ������F�n����ӱ����i	��.c�P�gq��M��Ջd��fݥ��5o��M��k�z�w��ʜ:�o����߰{
��f��}��5��	=Jؔ&�����7�d����k��J���:���wѠ�̴TM�ƈ����F�8c�M �2B����4�;xk�x@���8�tcs�J�䭺�}%�F��F���$4^a�=�f�]XfChp&Άk�ӂ
S�֝�A�Z)�?]��j��N���i��[�e\���c�qM���Ma- >�/�9��K�%"�� ����=�h8��z`�G�Y?WT����~�S�A.�7rSq8%]���*~v �#��;��fS$���y��j�d=�(�Ǩ�A�p��$K�s>)���}+q�̇!�
� ��_��N5��/��Cm��@`�e\S�x��R�r|���cX��p<�������. MVޥ���iP�1�:£���0��	�~�dm�����
x5���^�4���CM.n�'������1�y|KN<_"W�K�S��`��O4��%A������tX�tPr:`{�8(B�
�7��y$[�>
dX��-�Y-�[dG+��9�]�*Є�_P���,�g���J�V&�F����Jjx0����;�pj� �2��Ī��x�V��S��W�j�+���p��
>}�}�-(���U0g��҇��`�_,�V��{�3���ٔ�~��o��QR���B�����	���1����T4D�;}x����f���7�&OJ5�+�~�R	-��\��dT�����D������*�F��oQ����˹����\�%�@��Sj_岍O=�^�~��_�U�GR\��5F �E���D:��J��R߷��Mo�X\_Ճ��ok��(!\k&W_�J�:�+�*� ��b���O4��Jf+��G!4O�;�rN��o��f���S6'���rZ� C���}����ja�NB�}��f��{G%~�0�ִp1P���aL�������Q�� �����#4�S����*��ۥ�rG;n�.|�Ϙq�o�^��܎ C^|��|ł	~N�7��	$�S� ��a�:�}i�Kx��m���G(=ڂ3�ی���yw9��j5���/A[�#ALcE�O�*%zx�8M��xVT�F5;�L0��0>��O� �-�# AKTY��D�@�CN�}GX����0������$O��L�lg���F��x��w����pW�d�TS��kŎ1�K ��wP�dr<���t4�[��b[M�̕��w �U۵�)q���a?}[�Ô�B������C�~7��C��ާ���w�",��QUg��[���2����Z�[w?0�>,a>�����OЀ1�qj����U�]�K�s�ZgG~�Y;�CW��{z�λ���h%))��}�i咴�x�x�s�.��a��G`I��48�}�C3���N�lO4�a\� Ey��Ѻ�<Ub�w]�6�A�'X��A�� �ֽ^�B�s�-
`��Q�}�1�u)�\�:��u�/�v�p�A{~���K��8:F��Ui��$�6�6v��_�����3at]�UJ�G�;��-+"���y��9�8)S��D�5 �5��Mwlz������V}�y�*�����{�d]�D:@�l5�F����!�?�AF��9��qcc���H_Ѱ��Zϲ㥕{L��nv��"p-�7[�zPG��������I�P�����b�{�*�2�HI��r�iA���a��Q��4��W��&is�iً�O��Do�ӏ+��)#�@&���.��"R��!��&�Q�����A��	O�P"�i$�ux��}nM-I��S�89��i��\��8^Yq����.��Iwn^(}�� $z�\�'>'x!!�[q��'ʒu���hP՛��9mJ�5�ꯥP��NZ��a�ה��{ٕ��@���ϭW��;��0*Ƈ���Q�ҜGD�bb�C4�]������+b�C�*�;�#8����*wL{��/�
v.�k�.�."m5bK#��~�^P��|�#��L������������yY�0Еy`�I@֐ %\���r
n:�z�82H2 ;��OR�Ͽ�(����P��c�/Y0
�ݢ��GC����s�7�Rz]��ڮ&���dĳ蚕ås�e�T��5|���	�o�s�������Ri:���E�n=��>��n�8��0�� �+�������h����K�����`e�
�	z�P R�IP���J�^�S�!m�U��c2M�� ,@�&�;���HQ�?�n��y�Pߍ�z�9��PH�����ia�A,�Qit{_��|�)PB��M����7�X�Ă3~��N��:���0i��؂����,�|�+A#_����Yv�Q���C̮D�����SV��6ݑ�$8��cN��'�{+��/��yWۢ0�02̡�"�/|G�	߾�W)�Z�@ �-_�<Q�ع+_vv��}ڪH��z��Z}�����h���R���x��\N^��fM7F=�)�u᎟�{gH`?������XЩ�wt-u ��G�ml��o#���bp���݋틢{>WI�U~h���E���Jst�a��i��_@q[To�=u�Y��޹�!�4^��}��)�e��C�d��t 4�k�n�e� ���'pxS�Ū����b�ߢ���Zy-E���t�;1h�K���J��I��6�94��	�B�n�8x�vJ���}�T�eg��p���=�@�x5���L~�o��g���)�ʣ2`�=k����'�ϐ���Y�E�
��D��8w�X�'�g���<�
B� ��g���L��\����M�¸�����UE�k���t~�F���l%'�$1v��3{�
 ��~�/�u�$ʣ/�-g��{q˸A#y�@a��P.��������If`�4�l�ru ݭ�hO^o1�?a�w!�.e}0Й睻��&��,�ޢ?{�-*hB?/`<�Q��t���`���)��ů����ʹ..��!��}Eml #[:�O~�X�D'F���P={m���px{+�>AsL_�Nbo�W9���a%�D�\"�v�Mv8��rU���Q��YWkH1�e6*����D3yS����4�c�J"Ǚ������=��'Tۢgs�f��x%��z]�m���=	�wxJ�Ό��ڼW�H����
�(T�����}�\��
<���i2@�N"�:�c~��������j�=+h����Kʽ���# ����Rf{KSa%(G�Mq�Q�r���Df������u����+J/v��~��X�U͑$�g�����&-�*�6Y��៚p�<!��"�f��b�b�봕E�ƀ���Y2��6�A��������
�Ȏ)j��W7Z��%��u�-�!1�����G1r��lb�����֠�z�$9���TX������A[#��#�.�����+��(}Z�77 Zü�tLԁ�p�E�)#A4&�a��?|�J��ʻI_�3<��H�Ir��o٥���q���%F��-�fS��t ��r���M~2 m���sr����	��:k�������Ϝ�+6�TA:hFeX�R�%��	���tB�m�rE�	|ة�z�����t���K�#��Q̅�Z/ɡKV��K�r�0i�F�~��+���� ��_�ǀള@�,���/�º�#v���>N4�������!�MF�������+}�iF���B��	�pk$S"�ph�M>� ��-�ʯ!yD�a0���A��H���=��ֹ�I��o'g���ȳ��۝��s̢=kcia��g$`�i����$g��bC(<�gk�/J8��,�ת��c����u�MT-Pݷ+�tᤐj�^�7~�M󦬃�������ti�ҧ+��p�����+Q3�P�o��6�,|7��a�.���4Ӄ����� B��^e�6"9���igG���Y��>�L)%�h��I�k���,�w�۰�M$bi�_0���RI�y��-��)V�����MW(MZ��`7��J�����/�������u�����fh�y�Ů��L�)t��ii��^�jT���9 t��&�Q[���0�'�&�����͛��/9�vm=��,}猩.�ᬈ\�Ә�3am�����Fp	��Ene��A��[_g/���}�<^�z6�Q�RXk[M��(�R0� �#��Dw)�Y��t�@��IM.�>KZ�SfE`2�`%�2����2Zr��T񖑀�(��iQ؅�+�&&]7!�b�8����CmE���.`����_�lQ��soj7SU��_�zl�_�Y�E͏�������e*�4"�����.I����\�WD"������A�1��i���?T�p�o5t����f����v]-��H��@0�·����u��u�A��k	>��.��%�	�� 1[�~{���:��:������;�4kH�����E�%^X���D�5v��F���]8Ը����acӦ��	�_9��3J�uP� �B�+�
��[@�Q��e|�5k��ۯ�9.�U��E>�2*�D���Տ(�0�8a���yE�[���6��P^�Ҟ��y�K���Tj�#��|�([��/�	+���K{��@�]T*��?�8E�;�c��� ۝W�7R̃3���G�I��o�kpT�% ���8����߻MU�-o���7V�`lR���K!��"1JŘ)yoذ�	�
�?j�^=t�{{vKJ�����+�G�o�jZ���Sݚ�Za��#xK/ח�d���-�B�x(	��N59�dV����|��&��S�[-`f����t���8�k�M5Ə���E�A�-�� �.&8�˘\Q�C��s`���H�j���T#�'0�x	���)�2` C�x�1*�����u�����٠'W&�g���	u��(آ�J}�00&�Ƥ��癎��%~�em��*�@�7M�w�U�f*Ī|&��u[c�_b�{��:b���x2*�ʸd��ã-�F����*CYԶr��U	�,Zǵ�iG&��Hg}^2T�� I���Z�λ�&��R��%!�)��r��3h��;���1��O����C|�@�A�4�Z�?�~/�0�{��w%2����đ��I?m����g�5(�x��v��V��Qz� (��e��Y��tcF3%d4�A)�o۫�v�6)�4�W����DL��t�M"	1��s���l�kI��CcS�\KwB��g�}q�)��[�����~����e^�'�����G_%��`�uA�:>ܒ!0c����s��q��FG?�=�ҫ�J�����8ntd+��/9,ICv"�_��1(S��
�R���YK�-�4���l����Yk{��R���3%���8����&?u2�,�х����w��2��Y�l������2�r��+��Ĥ�U؋��'
P�,��N�n�aP�J�D���)��>߰i�����d�� �����r#�`�T K�ϭ���4�w�@���Z����/$�Ŝ
�|��eM���M�݊?�p����H��cui��舼��i`	%���rY}!�q�&)�C}�,"���W���/Պ<e.tXTp"x�����N��|�z'aqD)�����v�߻Տ�[�{J�e�(��"�l���B��ˎ�P�4����=�QQ� E��2�s5�'���ʣ�IOj�w�$�
�K{�L�����A<Oky�����S�"��n�nx��S���Z� =0Nl/70(�_����K�b$�����;�{�geT�l�%�٠ p�s\"������:�,>� �*W�*����qiDe �W�\�_�xʽB7�3��c���z��ҝO8J,�P��W��H��^��N�p�r��3��f-MO���D6,�����7@��wm[��[8g��K�q�Y���u����U�7��8�	�rK�ŌU��_�r)bj���Nf�"�$p�Y��,��N���)���:@���|$����a~z���LMڸ����F� u�Fԝ�(�"�7
�mn�;���DT�$��Ȑ �e�4�NC��:4����I$ ��z�WL*�9K��@��%�(�,p�t{�Y̛jog��'��@x8qPn5�1*n�)�6�Z+Ð�Uv���/�����<չ����qSV�E/���^�}��*����|A�Lj_�(��?Օ)$Pa��u�@�U�V�y�ۭ����9
��6�V�p��(g�>uf0E�����#�J?t�]�W��yᦡ锌��Ff���F#@a5���c^���Cy4�6��D�Bv��"�i
���e��,@�տ۱RS�G�������Zn ���%y-�f�_��:���J �(��_�θ�F��%�]K�!�4K-ZA����Ve+��$3�3�f���1d0��K0�}��v��+��"}��Y�w�Q�}.��m��#9˹9���R��ֳ�V0:c�5ƪ&P0�|���(�]m.�+�-��Y=-�ya�
(t�5DGP�\1ȓ荊T��(!� ��xO[��G�����a�9'��w�7�L�SVקb��2&����]�l���C5eࡻ�T�z�Ǖ��L��I4�Iٟ>�^��x���X�咯�l"Um,�<��b�U�˅~5,ϢuL�K4O,p!W�����0�c�Z}R��|3�\5��y{�O�@˒�%���8�,��X�*�zS�&�j�gvhH.�0��h9.��XN�7�	���f��;9�e'�tO#cߚ�Qi���)��ⷥ ^T5��F����բN_���WV5���.�'p�<3lRܟc��p���ǧ餍xsP6�����?����N<?O�ѻv$�Jț��.��}YP�Ҝ��{Ǵ��O�s��qO�����ĵ��ٻ�DBv�RM�W��A3+����l3D� �v*������ʊ�ÇiS-yy��c}��:��97�]e-�}���d��\�5)�S^�G26JvǗ��"�Se)z�r!˝��&o/B������5����
�d�u��m�����s�i���y�X��E9���
��QՕ[��X���yɹV�o: `cC/�����bJ|)h�=�?R_�L�B$����;J~zۉ	B�=C�D���ʭ&�2Ǳ@�z�?Β0ס���������Ѯ����X3�~��0�й7f�rx���A�إ=��%%<�|�t���w��d`�$|ds�|_�l���*#��+�~uMO�P�Vr�����Q�u���tFMxߗ��S$�����Ҁ۷���'@o%�m�xR��-�ӟ*
 h�c��.�,�����zゝ���Ok␠)P��(�o淁T��4�Pth� G;+ζ��P�,�'���6u4O�`T6z�A�tؕ�"@.�Ы�=�bř���y�jI�}�J�۞>H��X$��~n<N�n��~4�q##3�y�l�$�D����!��9'�zíHY
wp�����q�A-�nF�v�r�󌌗�ea�>?8�V�q�L����[���U?
�8ϼ��ESg�!d�JMe�L��JZ��	̣D!(�0	9�S�j���Ky����.�+�M{<����*Af+�o�����e�6��,�bD3~҄Ӥ��,���%'�$�q�[���K������h-4&�Dg����������Ӑd�&=����Qip��F�-5�F$�g�:�X�lC*#��L)�-ј�����&�WtSB{� ������_�<�*M{��&d��i��«Ce� Ǉ
r%J��(-gz��Z$��ဲviI��-8��F i>x�-2����Y⨾����M�[�ѵ�r�p�qt���Ę..�7K��[��=z Qp��A��3���c+N���'�����9	��<k���{�k]���;�x���Cs^��������2�O�f#����	�C�a��C�����s�[o8>�{�DD��ԾX[��/��62�a������Z0��#B#��=�`}#��'�������{T���j
�!��Z�5h,S���Ǎ��\���f�c�i�����47���'�����s��,ᵥ�V�|sz��}�p����P�/Ҳd:�;䭓|�$�%9/[GbFJ�r�z��=����(�TIHw;z�\����´�f����͐U��B�3,9k�){�H����wS�����xe��.�\b�R@%4C��� �wh����iJ����9,D ���Vu�+&�-�@k�x�����-�>I�%�}��m�p��ob�)N�������jR�镒��sd�d(����d�M���lD�^C��5�,<��=ײ�6��&���>�¯%_�:���}���� d��N?�]��5��]��2KlJ���X�
+�
���:Nڂ���`c~������t-���Ш>��Q,OK�9�Q�|~vת��h���T�/��GK٦�ʰ����;�v*��t�M�����>'�Ib��ףT11��-	%�e4��>8)z�E �JÐ[k�,�q��Z�3
{ ��`���F-�E��=��턄$���Q��g���nA�������)`+�?�
������nK���8�1��;.���l�qB4�nαq�B��c�)f�ԠRcK��$���,���ǀ�8�fB\��P��O�}��q�KF��B-��.q����Yt.*�_���AO���,^"|[&p1w����\y�����It�$QC�m�����������Ґj|&�O�tO�Kv�+�M��`�X{5Z#iIkx2G�����Q1����?Ds$"�@����1��:�0X�����K`�E?&��SAu��ƕ�"��n�!� �1.���aI�=��j���ۂN-o�П�����0�I$U4��*����.�)h�	��Y�g���q�ڱ�� x��=�
Ģr�GW^:�s-|ҝ��'���1:����*�I��>�}.%��*q��N�o��|��U�����^�0�/�oi�}��!���٨������_v��zJ�Z����f�,���Q�(v�//O+��2N4��ɞX�'��i�,�3�6�q�ȿVr��J?l}�޽��=�+NçV�<�W�����T��I�Sc�l�Ӗ"��&�F��6w��]K���>��~1�s��hP����[#�ϱ*߳�x��XB,6��*Z}`��#˯��H�3�}c��_�� �_��۸�Fs�;���E@�&	��_�� B��tWk��2���{ۆ�����q�9����ҸU��|.�<�m��ax�*u��e�v)�@_B��?^�Bd����~d�'�6���x��������ci�3/L�"�AX��Ѡ)�&�P�?��u��+����1e�N�~q� ��{�d^����
nĐ~m�	�������G"?� ��f��V��� �K������w`a��3�	�$w�88]o��,R��zk�4��׵?�oG��/^V�)]��;` ���s�GĒu�MW	��y㮾d�x&���~kC_^K�G �Zܚ��,[x+���S�ՂU ��q�b��M���@��z��z�S��cs�)(��O����!L����M˞?͆m��Q�� �񛚲��c�
��������_���(,�6����eH��
I��#�˙?����',<Y�e#���:��K~�*TIPEKo7|w{Q���>�ˊQ�t��(Y�kҦady@my�E%�ܐ� r���M�3*&� dqд�H��`�ycύg�Ca�g���:K,�qJ�5"�=W��� ڻ=�����PX9A��Q��J���x���Ah�@2�,�Ɍ�����{��8�9��&��&u�UV�D��
FZz���f
$ƒ��;V;�Hb�K�hme����8�V�������s���0�7c�Ta_p1�e��$�������"s�S�bs9�����<��O��fѬ;$�|Tm�>�Y7�Xr��m����+usʍG}�bMM�g9�y�L�׉��qo}�zD��8~һ��L�
���tU��� ���SL3wꔨ��7�M��Ɨ�g���z'k*�1���J��[%�Fz�WP_$� ���͠?-BF\M�1� k�@lW�Ep���jg7��8�sB��/��$.�O�H�I4U"�Ut�u��j�A^}��ěMS�l���Z�e��VJ�
�O
��.3eP��� +�o�񨖱y�{AX��L;S��U�Lڍ��FH����G.��ـ�G+l�㕷^ؔ����ҥ(욏@�kH��,W	���+PYX��P��y�(tL�'��Е����v�^����H����2�*g�n��Z+�t�a^d���b'_(c�Y�Vu i@|���۾�m�yT�Yr�K'�D��k�[LD�XR���	�D���(d��aY#��"ǄK�C����H>2�?��Ca������}��?�o�),�0n��p�l:u�Q��y�
� o�ORg��h��9FUA2���r�Y�Y,yx���..�빬 ���i�`�3��1��DAD��BP,x�����շԘ;� ���)Z�pi�:������Y�h�,9�j!b��?��}��T_��J�3���M�)�1WhEe5Դg����矖lG��'Z	��mL[=�g�>�(|��z}����/l�W��lϽ���5�`���Q�+�Ս^'_�J�Z������e!��v5$/�MF*ՔF��Ԍ*�Bd��c����U����|����z�S
������"0��"�z����s���|�"����r��<���}�[��>k%�*��p1�e6a�ǹ��Bs��U-���<�d���]��x���Pw.����K뾖�:5���\0��սb��-mYM����)I���E�c��w#i:� �I0H�Y�g=��vs�(N��a������F��h*F�9F�8L~�YC��ٹ�@��h��+M�G��Ţ>1�ԚX���IV��t�:f�iܶߊؖITZc����Z,�q��J�M�O,:�
���v�gm��O#�Ow*;���I�7G�P���Ѫ���/��;�be�CFJ\�:�Qu?I�s�/��IG��Q�&Ǉ7�i�i��ߥ	���)X�-�MG4�$K�|`��M�nڞ0b?~Of�@ˈlD�}r�ټ��'rl{[��R^�R����ٝ��~�hN��UD	�j(9�j��I^	��8���+cG�b�����1�e�j�Ԡa�� V/.݋.��?���׹yj�Xd��!0T�(�c{����]j�wP�GvA��Eͮ����¶֮~y��"T��`O�f����h�N�`�X��T��h��M"$��G��~�f�!�~�S)Ѥk8�8����\$�-���b}�uzyB��Ut�,Mf��/�S�W����o�G�2�˚��� B��k5����wTN.�"M瑏6��	����'���xd0#���X�=Cy�f0[S���%�Ⱥ�E�Ja�0I�dP�7l��ƌݻJ�s�n.
� �F�-x�<�9kr1�棏.o� u��N p>�h��i��ڜ�Y��y/�b�O1+ԥ�R���I��N�	-u=3ɓ���Z���U���$�iL� hyI�Cx8rW��[	�v�x�k������5����6��6�Y��c^�� �Ò!ы7���H�Z�T9�\��#NTzjc?ڭz����@��͜�cG]�a��x#�u�^�ײ��Dytu�T��?NՒ>Lm��W��MW4�m*��n`����`<��3�S�GY���$��sA(��}���Ŋ#�[B��Q<{]�V$���q���� �V�LM�s�.� �YJ@��$�*znV�1B�y�#�B��b�W��Lg��!�(l�b3銡Xt������􅊤ã��;z2��sV���A4���ɳ�Iهk���.4��}k��I.08���;�,�q\�W3�pWQ�	^6�h~V?0�7�c�Ҵ%��E��"1G+?�i�"?1vI{V���y��i�����/�{�,I�\�-�|�P ���E"��+!�z{��0���v4qE%�Iy�?++BȰ�ZG(�l�7j���2NL�I ���(���R�����e�){�S=����^�#4�y�>��p��u�ٵ�H.TE�А��� �'C�_pܨB����A��Y`�`8�8c�QL�|@�&ק��Ɵ"*���<Tў����;Yvcw�O�O�0��1&i��#�P�N��qԦ�)�S+>U9C��U���Lk�K�Q>=z�J��I��͗��:wIP0qO��b6e�u�Lv������k��/q$~�>�;�p�(8AS� 7-o����!�e���O�c3.�*�l�G��"a���632�c��|���;�Q7���L&�H��b._��*�`GF�. �o�3mo �h&��#��u��7��Q���T�Ӣ�����G�k������7�dK���OD���:�}1�ڂ�p�у�4��'��<�/�&�Tk��
߁�� �ҋqAF��.��;w��~Hֶ�==)۪~3����7-�Zp��^���Q^-Nb�/����I�yC�VI)��ys��4�i��#��! ��+H3���\�,�P�ͅ�%[g�85)������ԣ������2�у�0��=���f�kU�{[n0��?�+����i��n@�ጮ��@��k����w!�?�7�@鹂Ӓ>ix��5�i���H~1�Z�>��ŕ�^s�6�t��>�C,!�@xͽ"{�&E%i�+���'����<��V�^��}��s�%B���M��u�&�V���������]?�B����/6�KTm��~��-t�����q��!6��$7U� Ǚ��gk��ڰb��� �,���s:݃�k�e3����(%��m�p��c���9}	��0��*�̩���m���"	�Tt����R�L/_�HH=xJ����cM��	�1�_�6�B}����<����+>ۗ��:1QV�S��H�L������n�I�Q����ޢ�� s�g:� �4SM�r�	+gr(k��V��8�7I� ��RX�xf�+<��g�	�1a�]˩V܃�_�q���	>��b;�A�'���@l�g����Vݥ��vO�W��~~�������x�?h%({��e}�-���DMF�*o����:��J�� 2��Im�V������'lΈ��,ݎIF�✧Rvt	�7E��77�S�w���U������M�:������j��B!�o����BE4Ye���5��A=ł��p5�!i��v �
���N��K��PP�'_jh
º����<s���lan�5�ȡ�Ҥ0EAY֑� ��Kid�;.�=m�����ժÞ�i�5�9���ك*��@�s�3i�c�%���q� ��U�#>4~�� � g䣫Qy��� ��)?t�?ޖTO�ܤkpGy�E�"���>1�"���í�r���� �;8���I����2�ɑ�+?���;];�8R��z�]���&E�ٮqA�T]�#$�R%?�aR �����, ���w�F��V��J!�{馋�W�z�~�ZGg�����n�	�0m�%� ~��Q��_6|�"_622{��	�m������-�<C�V
)�s���y��ϝ�`��|��7���o�d��I^a��aۅ�Č��t������a���o�Ě��'� If��=�}}��逰��E�%�4��i��u-�JW�2G	X�W����F�QXfr�"So?%%��PNT7���_n�KV�vV~j}��A�E��S�g�7KX����V�i�gU;-t w'�������}�M!b�4Y�I�VK�׳WD;sb�e1���o[��p�ud���͑�q.Q�"7�$1��r�P���>�q�_'�Iטr�-uhN(��| ��ާ[��jff]�� ��"�ZbC"����ˣ`��c x�G����x�����g�߃I��5B]8��@T�K	m��0���Q L�_C���qz*t{��7�߷�FR:m��o��9�����\�Zx���\�:�\]����0�r�4/�j�q�#v���8e)����!�֕���2���ϒZ
���l��܀�_>��I��hf��ꍧVm�?�_ 9}QBGti��#
��M$U���L@��ҁ��2ӗz����u��m7Ҿ�q����C[�kCb#rm�l�#o���X\�%L^d!|K��[5/�oTM
���h(8����[O��'�y�F�%�z�2>*Kh�Rҽ�6���k�pV�@��l���4�z�4���$���6<��:�V�Ϸ|����'�^��}��K��bK{x7�t����c�W E��1w�>�Y��u��w��ESU��
�c;�7
͓�ɣ�֎�A[�����e����1ha��ܷ�����=5�Y��R��4y-����v�C�V�"��;�fn�,���r���������$��9���z�լ�~��Y�����5�p�~R�{Z&�e�OxXOe�f,34�q�'36>D��ё�"	BRq�M:pPtal@Su���ʲ|�i�&��F��L���J�G&�DG���.��)iI�Hf���@��`�\9B��8̭�
��c*-R� �s�xD�v����a=��:�{
	5|v�-����ı�������sh�I�'�U���]q�\�;��L�n�:.�������%P��[LuV~Pu�����o��"{������n��^��66�Y[�$�).E���,��ͨqa�|p�;�Q:����1󓡴�ʧ2�Ot%�}C2��Q���6�(�m��9���\��|'����K�^�Mr�7w==t�d]<W�A+�k�	1�BO�VWMn[��3�󙥪�Gm���MX�'=5`N�z�n#J�*��>�=:��y'#= cw�F��p�p��Q��"g��W���@9�p����܂�	B6�D �ӆ�Q0r0��Z�	 |<�I7}� *�X=��U�$s8Rݞө�<Z�4�/�d+�L��j��S��br��v��c��^j�!8w��Ax2W~���F�|,�7h'&� �B�ԋKn����!���nx����fe�QN|P�|r��:�=�2�w�9OxW3��CF�xX_�h��~�IU�����#�?VXTWW�l����ݵ��/�>Ց��r�Z ,���^��kv)�S��W��I�����,��E���i�I�N�X�a������Bm¹SH�|�a����T�cq����o�P&P+�-ș�../��� @�G�Ŧ�KKҀs\3?������n�@��6�6��	�Ti�����l������Uz�(T��
���:T��27Vƾ�� ��qjt�xb��Sc=���%VƎ���P+�;~�0}����-ӱ��U�^��ѐ�A'����XDJ���w`���%w�F�A���l��҉U`<Ԃ�L�����v\�f���R#�Be��]]d�h�f ��|E�2Z:--5����/�;fbt�������YH�@qѩ�Jd�D����j�	�)�
 Slt���Ȉ���jL9@�5�����p�5���r�Rb����ᘝ�N1�n���q��ջ2�'D��	б�HP2�"e��c�|/���vK���%�9E�8
�l_�S?Ť�?ٔ�����F���!����l��wd� l�w�.�I��\��@�y���=2���ġ�;�~=���D�l��cr
ψ!3H(N@;�{�iv���vb�6����5:V�7a�ݻm���7ڶ%"}�:$@��e���\8w04u����r�|,\\����J�*l�@��n���X�jF֨����b�����T [|�dO9�}�#������u+.���NTQ�{f�tS�5�#2�I���B�z8�ԛ�oߡI���/�x+V�w��`I�KOODݹ�{2�B;r+�ö��R�x�)M�$�����#�K���'u���[�b$��M^��E�ɻ���F X� ��W����u���H�˦:�z�F{��\@8�bH�*���%��[��*��c9�$��[2�?(�c�䂶�<)�;��/��&4�m��#i��
�!Ų~k�'}yEb*�fJѝv���Dc忘���t���0 �NicW�m(�����o!����!1�_$'�ޞ2w���О��Ŀ��!�nb��c�4�]��/����_w��pP!i��>&���M��/aj�Z�7͜i���mPkrK���T������Μ�ȕ)Ʉz2L����装s\&Ow�:Lޯ�7:�L���G;���t(ğ�)@����{X4F�yT< !�9?�j`�_��L�8�z����l�H�����T�eHT�C�9��W�%�HK�?x�぀GiHV`~�����T�m�G'~\�������ٿk����r��L���]�y����]� @��-:�-Tl�O:��<��~q�J���"&���`�5=\�p3RF.����F
�F����n�	��K`C6���sm>�H�(ݐ����]zN�\P_�8;$�L������e<�����t%g)������V�Y��b?���c�~��L\�	�9��3J�OaL���n�9�;�vn���'�e!U��%�F�B�@�Nb����Qn�F��pih-������b-�/�l��~t�?�ĥ��|���
�Į��N�[z+���p� *%��]*C�ӻA��H�ؒ��}����\��|�b<�G���oОc���qt���X|�[�@+��l�'��
�eڐUO����0*m����3��lLLm�浿�mЂ��=P�r��D&!�Q�up�2��	�X��a,���`�@W���]���ݽ�R���*�Զ2����L���7��
G폳P�L���H�(�nCgj��}|Y�&�c/S�m tT�V��M����W�ħ����D��[E+��@{��!C.]��O��謳�`
��|���h�ZC���� q���N�r7QEX�{l�Xܖh0 �J]����C2W���":��D��jpӖa�+��m�u��+}�IG��re��TxaD�����@e9u���KW���>~v�P��i+��M�J�'��2��@-�"���_�*-K"��J0�r*�����.��"�v�oz^ԯL{�)�g1a�`{?��7e�:O�t�V����_߉졙���.vWAx�/��\�WH�m���<�9[��n�������=��Vo-U�ǥ�M��h,<��˖ea��	���D��b�&ȉ�����r���\5
ms�+74�܆�2��9c�^M��D�����y(����r/4J�*���6ԟ#�Tʘ�Ý�Z�w����gv����<Ą�+&I_ȭ��h�FcG���[GM'���a���O� �z��SH�}iM�ޘ|F�F!��	*rDi�gn��[�𢘢~�J���q����UyYZOCV�'4g{E6bI�n	���J7���cXv��Z#�g�dX�vX��V�`c8��("�2J�x<���Che�n��c���C[��]۴A��[�G�C��]ʾ������*��5C�,3B9�.��u��^8wL�3�����#m����oY0�E���Q�+\Ǖ鶎V�IŖ��j�1�P�1���J���!lЋ"FH����]��u����������!I���"���_5/1\��>͇朣��a���Mf�X�_}��5ćN_p���K�b��$Yo��(��/��q>��]��������>/%�*��󁎯�ɶ�'��-\~	Q�Jrr��t��n����I�;&ӗ>W�P,)�8\�{ė4�$���!b�°�<.B�R�Dː��%j�צ���M�+>(�֖4d^�z��k�Py�C��y�A�,��݇�I)��|`3%j�O��S�0�L��g���i�xsNe;*�VD"��˧���)L��Ĉ��%^\35����X�	��4T�Mf�i 5H�t#+5�s`�C�����O"�ӈb����B�b����K��Rs�,Ӻ��	M�%G�=�]��"�e]��o�kY�4��� 2��6�↭��_�klS�nB�/dpX	D��G˚����x�����+�B?Y������l��`3ɱ�Z��c������UD����޴�@[W���h#����=���ڑo(������D�) 1)��i��G(�D�"wê�&`�b�Nk�o9djr��V���/��a����6y=�����ܜ֦F�X�MהsA�@�[�6ׁ�xh#j�3�N	��(���Q�ܸ#�R4u}ߢȳ3Ö �uP����,۳Ѫ�m��Ǩ_;-�&?�jS�����UZ�O����,Z�jo�	���ʕa1�Ď~�'��8��������C%����!<[���kpէ	Gb�_�_���S]`��bP��N�{�q�n&��_��8�|�U�ôj��\��?h�߃g�!7��.Ǜ��<O0.?=�r����Tτ@+鰐l�YA�"o�]�|��GI����Í#2��ň�'|~�4o�}�x��6ܝ�#��#^�z�O+�J�d_w�V��(�O=�BJ�&�CA���UR�njA|�ʗ�pk8�K��(!�;�Q����Kb�r���M��0 ހ6�����!����,��J�u������i[�����"�-	J)d9��/c��P��Jq���Jӄ�>	dng��g��QB�@��}�A�4���:#]��s�����/D���ggu��û���+/>(ᶦS�����rw����TϋCq���@�r��*n���iӵ�����I!��#"�O�+���p��6����7�`&���kd���o�_�p�>&+7��Ǧ?<Ҷ�2%��=%j4�	�l��N�-�`�|�y�m�E�M���a&	$�)�����(&	0/���j�g��E�7����ӆŷG�M�� eJ��vZ�
��� �kG]5�*?�]x
*%߷�w�mt��J�?���*��b���$Q=�Z��1
O@\�dg��_l�4V@��ē�q޶�l�͋E�t:~��g�e<�ux�S:�,K|�u�,��-/c�mmu��54�<�k�_LU���y�@k9��G~��8�:��%YO��LG����+��,2�,$JE��0�5���Q,�_��@�� ��]����:�; �a2��WLZI�3
��$2��}�4��%%? 
��7#c-��r���o���n��0*w��1��5��mXR$@5-_��b�&Z�Y�q؇��R�V���2��N��OK[ݎֲ��3<�s�+mY6��d��V�ː��7|@�Z�B0��r<�OA	0%b����￐q��x��x�����pZ�-���G���e]u��\�7�.��;�"�u[�cFv�6�Q�|�n�&*(���G6��B�6�lj3�a}亿�h��x�t�A�	oº7/ ����j���b84Z��0��(߮�5q�"�#I!u�L��nJ3YU~ae�(�K�i�������%�UD٠M��9��<��n�/�܋e�|TX<��P��b��-�OS�L]��π`u:��:�����8�/	��1�C�Q/�PT��E `�����TV�{�E����es
��X�h���[`����61#r6�;~��x �9�����Y�2C��u�vd�i�)'�ȋBQ�@qӶ֧������/K-s���f�"��2�"
��6��C�){��E&^�ik���\����F����C��������|kP��y�}�5�o��Xz6yx3������BV�vQj����f����`N��N�#:֛nQ� @�����~i�c�������X�� ����E6�ޝof��9�p��x�N�?g���2Y`��A�V=��ǀ�/T�ܑ��4ד��uպ��G�ϧ|��F�U���j@!��&���ⵤ��5LE�_Yw�[.KS������/��5�OK\g(��5��g�E�F\�9q��p��Ij����)R�g.S{֋
�co��bMy�/���|"�ű���iA&"�d��'�j��6_×h�ڦ�8�I��96uo�m�����f��x߾��fհ���!��ɑ�Q2.;�� "1+ +5<��0
*4�<���ɀW���F6N��7�6e���گj�Y���3��`CQ]�x�J����1�_��������G5���;��"Qd�
O��z���?�}/BDA~�sv3��G!Ɏ�r�%��2Y��-i/.٘��ᩰ�򅭓��6[��Z�Џ;3Z�L�*z��%ȥ�m؃P6@��4�8|Arc>������1��vz���؞T���s�������A�q�[9ߥZ�{�}+�%K�G�WoE#_�|LO�bs��*���$�;����~�d�r	�Sý��)����Q42�$V�o)~�����uĊ%^�n�U�H)1{���j� �����D}T��W�D;Q��	�4�&����k�/A��ϊO��,�̀VƵ�mmx�u_�x��ґh%,���{�N<4߹�Ӭ �{$�a#au�E6u4��[��IcS��K����K1�d��`�{��S�?�l�i=��(�{,�|�� ϣ�o��G���B|��Yު>	
s���8��g�Om={�{��|֤J�=�	_����T�I��ǿcزzc��i]�\P�j��Gv������Z���t�D3���	�Z1G'�7ud�7����sɱ�f�o@�9��m�y����t�?Zp�"�=z7�(�"�_�Q���H��1�
�������)(�P�� �.%�п&�BXs��¹�/TI�z?�I����E�)f1������-k�D��������;��,���O)�AD�R.L."[�C�1�d�j�v�	¢�0۰o\�ҌY���:=��T�������p`U����?\pI�W�4��/wHq#x�/�oľ����?L����-FYڱ@bA �)�1��5�~��HWe(�$�n�U�<֣��ZEZ�'�VL]��AEs�:B�0K�43�R�_Z߲E��h�\��m���.0shzX�P5���Qx1��r3�W	@�~2��}����z���'O=�ɬ,�?d>X�SDS�v��/Kٴ�wQ]^ϔ]�#�oT	2ڬ}t��Ǣ��H)7~'�1�2<ZH�&���n�:J���hà �|�W[�R��i�读�y�2��ٗ���١�m�'�t��~H0D0�.����28N{��3%Ā��~��*V��r�	T�j3^�����������D�q�+j�ȡ43�oo����xii@[]���;�Z�����`�P3���r'M.�ݓ�8l�xq��/8E���@��h�7Jl��+t�ȿ�������,)� �O��*b&d�_=#��ӓ�.����p��/�6ɧ`��������j2B8�q��tM'���|�i�ʮ��y�N�g�[�6��I$������Ё�Y���&D<whs�����	?ax��-
��(pΝ.G���x�P�(nP���sNɶ�\�(s�ē�P��Z��dv5I�:R�O�}s�l�z�l
h!o����S�ȵ�b�qh�LGT ��U��(W��{-�(��q5���LS���&��C������g�&����s�|�t�+���.�d叨�C��XP㇗��m��:ziK� ����2r�4�
 �+1�Z2��]�h�̀[�y�SA�?�2iu*�k	>)
 # �~6R���ׇ+���ͅ�<�I�ӊ�]̮���ٛs112��u&�MQf�s��Q
�/�`�,���
s�dc���y&�]c�at��f*�;;���Gm�V�ɦ�,-�-������=(f��NE�V̙��;���|�K�.�̆����h�������U��P�J����+W��7��CP����fBP'����/s~��$l�1*�-B�a�s�S�]=�QZT�1���%��#�{?��w�NP I�(�8�ʖ���$��"����/��DC��Үy�^ᵊ���2�7��>�X����h�MӴ��0=W��1Pч�=�$���L��N�ʥ��Q�{1Y��@V�h \��y�f�^T���A�3��~[Z	��Jٜ*l�5<2��������H�%�KY�Pr͜SJ<�;ZM`m>���E�݊�#�ro�T4\��vt�j�V�]|U��cAr���kz^8X��b+��|7ڿ�t1vaN ��t|g]	�N�*����q	�{�\� �nf
4)Iq�{A���?5��5]Z�/������
��a�[��ݗh\�d,� �����K��0�MâTB�,C7"V՚n��
�)zy��I[g�w�~@��P���-|�d@S��X�v��s�9��*f��`H������.S�%ܜ��S�dt4'][mC�<L�]�?�{�1o�#�\ŝCjM�@�K&�+��@Y������n6�����P��h�YI�#����)�ܳ<g�w�+0�]g��!	�Q�8"���ǩ����1%�c2iq����>� :c�)c	�~yȰj-�k͘n�Ja����5]WZ�E�ߤ�n��n�W�2R�Dn���Dk��}�(�!������M�.�/j��*j݇F���YI�3)<��/��~	�'fA%/@r�{�㯹��&ދ�q�|�V^8�? ٣�w�X�Q;��U!��>fX{�����������^|��F>�hG0�)��	(8�j*8?_�����L��kljRS?ƛ� �Ie��m�rs���V� ��4B�I�r?��i�����7�q�0���:��C�c��C��31����T@aL�T���2E���+_���#R*{	�nUs^�$��r!�\�I��q"+����')ZBs�bWh<�-c�'mO6D�Ro	c�)�@l��|4�On
�h��yE�N^�3�w�<�%&� ��J7O���,��-�2�����~$�w�4���\�Q^�ڄ��iӂ�0�y�%^9�𩬥]�20��D��������dI���N��uo�D�)،+��,��e�IŜh��V�x@��;h��6��:�P�a�56�[�ȩP}�+�����7�A�Id1]��ַ��%�Wc硟ju_�Q�h�mW�~Q�����-����@���V����p^%YD��;��y�aY���|����7Y�}��yL�ch�(
���1gm��G�%[iA�*eǳ����-�DoN�,#E�}�e\�������V�)�b	�a%�FF�k��*�'��f��s����$_p4�d`
����n��Ar��g��)�O3�U���l��}m�H�U�f�`�+��	��]Y�%4|�+�! �(C({���5Mp_y��̼�rݔ�p�����M�1���"S���U`��]^�Wgz�a�f{��-m���HV�P:�K#��x�/�/i޵h���+���B4m�������=��Ex�g�����H��6z��@�j�AmĚX�!�JP�g���u�f��,~L�Ӱ�kV�������|�~�;�?���-ּ����ݏ~��#�Q�������V��m�f�Ͼ뽧'N�����P���h	��$�>	Q�7�t=����Jօ�!4��H���a�!*��n]���[�r�Nf�z��ZXQǐ�gS��5@>zJ�$�W��|���8Q�(7#�۶���A~QF6��M�V�=�ޗ"�%D2��䧝"��S�
=���kF�9%���L@dZ����H���>a�p����i���]���u���E���
E���K��3����gɳxȴ��:{ӭ�ir�cC���qz !��X��s�Do�4ق��ZO@�k��]��z�)�p����h>w�

�@"r&�XG�E�ӳ>������ � 5!ǡ��=s�#-���|6�y�}���UyCy��P�'y�&L�N���
n:U����{��i���8E��E�N�K\[LViR�4��G�.�tV�4١�f��߁|3�۴̪C~�v��HrOvRІPi�$6v������|L�K^*e�Ʈ���tT�u�Bc��f�9�G}%�(�y9jN�vV�1¸P Up4�#�j ]H�U|�\�\[AJ��C�g�z���R?<�B��+�0�\;w���7W����;�F"� /�Q����#����L�vu}�y$q��ykӏf�ҔZ�,R���dc���v;�H�X���ã�i}�^JW��ﶏ��Ӌ(�9���);!R$��n�W�ru�b��MD�m�\@r#ze*<���!��e�p���͔)&\��vU%���ma!����,�J�P�#�%�!��HP�1E���W	$�`z����V�4��*��T�x��jM� ���0� ��j���i���Š�쳃��%�k�.�����'߬��s��)�?"�_��Ҭ�?QI�5�e����!�D�Q5�i]��
P����{���&��o	i�yZ��B�_��QN����5�����L����Z��v�����Ǫ�7��5=]O�����������x]���ش��ׂb�̏�}���Y���
�\�0�F�H8t����}�,�~{6E�=��Hf��>'(��-1�QV�\�,Zhv_��~�X[h�E���Ꜩ˨�?��xv:i4�c��Da��%<V\�(�ԥ��T�%�����ޤ���*�\��UU?�d�^�]�i��=��o!�<p�H�� #��sd�q�������h� /o��d"{�;۳�4v����#/�ٞRܲ��K�D���]�g�^�� pd��U�Nk�{	�,kk	�Z�:��rq�5t�����1+���rhvx�q.��"!#���������i���� �qŊXи&����b�)#q�0 �d�U*���t"����Ԁ�U��$G7�����&������ؙ��PG@g5�±������!+�������(���!ߋ$�u��60���>!��D|�j����F�b�Γ��6M=��J���B�Ì+#�)�t?�|���d�����d��=x'y���u$�����g���&ݹ�9����ڹ��>]k�������8�p��w O�Gm_�����EG�k�#W�vh���^���1�1����u��ǯnP��~9��R"�5*X��4�<�M��C`�����p�d^��b�>1��Jty�!j����N�����\�B���t�����6L��v*3�-�LFVVN�V�d������Y/����\�j5܅!O,����k1����;�8�c�2�n�7W�x:x�20r�փ���T�dx�Z���&j���!�r&��Ő�j�t��u���c�������Nޘ&�亸Sq�0"��O�7U+F�AMD�c�D
�X�WsAwWn�S��K���nB�|���W򍰁<\�N�|g�<��}�o��1jC�3*�dh����R��{~��Sz���:ZONc����*��O���/�颸M���h)[X�ԙ\�C�!Z�Y����68�ѻ�5�]O�s�^R���K�iS��E5� ��ۆ�)m�)Ќ�Ć;�CK1g�I��5}��1V~x}s
�f� ���fy`BT���f{�IɁ�=�4V5	����}�n�����z[�E������p�ױ�'�gA-R�u1ʴ[
�CgG�������h�Jf.62�-_t�dfT�[Z��W�,�s�oS�=�PE��c�HML��B5�!�>�Kv�y�ªq{���]�
�(e��U� «Ag_e�<k�_�Y@9Q��I�����H�ka;wl��gLK�Δ�3� �׃ q�b� b�J�^	��h�d&�2��˲S.GU��>��s���8b��KS�䍀n�.1s�`�!!/�,����G#���Cޥ$�v����N4�ZG��To q~����_n�nsD��3��%�B]j�!D�V������3�2ʹB�Vw�1�/Iƫ��vSe��:K�1���[�P_d��
O'S�-�.���l��*B��r��^E�>�CBs�s�N������B�&�Xe�g�Lq!���Ò: �ˎVd�U�ţ��U)|��qK�m��*�#����K����ֹiE���`@<re�m��^g�|���^a�����w�$M>c���
ze���;/d���T$��g#`���	��"�%��8�U��fN�:M@R]�!<	�%�1��^�x�w��N��b�Qıl���M9�)4|GŘ�����DF�a$JN�$שn7�|p8Բ,�뙝 �1�W�v�-ｂ�����)��T���nu8`pd��ڋ�=L4ޯU��qIU�̙��G�h+!н]��Vŧ/����9q_� �L8�m��_�OH��ܽ3��F@��A3V��w+������n�/��ߨfW5 p��iʠ"n%kR���'�a�s>�5u�j�i�����Dc��y�ѿt�J�t��:1Y�Bc�~go^ �>�x���p
�X@XϹ�{���4�>'�Su^)Ջ�U^�*�����q��ƻ�洉Wɏ�*�I��RG3���.$��dG��Q���^
���x�	�Á'���}|��>�M�ν�_�j��#z{�)�;�[u�G�^��
-�l!>��.�] ����*f�}���+ӲS���J�_�T�M�Hн�hw���Ե�L?ђ�Y���G,��Z�4�A%�,�;��?$��!�9w���:��^J{�t޽�x�{`�Y_v���|2v����,S�=�T?(�0ej�����5�1����\��+�o� ��V�#�g�+V���X�<X�H���p�Ƕ"�I�Ǒ0y�*��U�p�7
g��6�SK��7!HN������B�f(�
�xG�����
�-�!ʝ�l��Z�я!Ī���0Mr)�ޱ�|����0���13+�]ޠ��� $��{z�ߊ7�p#�cb�����Ь,o��=^i:K�o$���7�z��b��ٱ�R�Ŵ��]���/�Ξ3��/�v��x�^����-���sE���ZKf�#��8��ퟐݺ� ��J�\2֍�`���'~u0�]�����$���7�p"/�|��yS�N��Jݥ��n��';��э�k�9�h�]��ڻSs{��Y�;�K�`�2w�㔱�U�=�р��	�Bn졏%c1��A���o���� �&U�:����&_�
��:	F�S��
BY������6	^�h��N�ϧ�(9rBH��Xf�눰�:� �/8%�j�1�-� ���&(�káD1�j��6`�i!�ͭ�U�DO~��2~F��N�H�˰���MS��9p�S��eM�Kq��ے�!�È� �;%���S���b�^Ӛ��}C-�Um��[U����y䨋/Ҭ��V��RW�<4m=?�Fr���))�� ڼYZ-�I�='��:r�<��5I�K��@،������bM�;F'�B��'�F[�M��7K?����<k��_v/�.-yL�|��(�T��l��C��)J=m���zQ��d=��C!j}���f�B�)>J/�6 ���O�ˀ�w��c%�7}��G�_�2�7�4���)����_�9�W;����'pk5F�D�����X(��0oM1�]�j��(�ޯ<�[�ӡ1���;� `)_(@�-v�^#릻�P�#�8�����		U�לhI��q�D����~?��)�G!�~��bP��I#d֎X��#Y� �⸔x��B�\$�7"NZw>��Z��A$E1n3_��n�����N�U~$j �5[b�@��O-{��/|n��A�ꈠφ��=b��}�-	:�%s���2N/��D�q�N�a�l]�{��GK�^~����H����x̳J^�5�_�w�PP|�S95�1%�+xiچ��x,,����z�R����;ޢ6��2�C�`/��I)bۿ%v�Z��df���>�Rq�!n�����㵯����7��BYm�o�yrB�*��V�EV�잁��ƻO�3z�q��ߒ�-		���s�뤜M^EAY�pj�7>�[o=k�w�����Y�k�K�R\r�ҷ���ȗ���,y�Ex7T��I�~�
2V�(�Lڑ}X,�k�\��<�8�`���N;���jo(R���A��+�#��!A��P�+)0�X�M�Hl�g^�x�62[�Œ�*'�;�6�p���8�!����tt��	�W�i���k������ZK#|�[ɝ��Ҽob5zջ�
���7�j�]���q�d��Ad�����F]l,�1��57q���=.�sÂ�O��T��g�Դ�O{�vDs�oC�X��Iy��_�b�M >%򫱹0�� �1߂�RQK��R�j9c���7V��_qk����� 
�����>��f�}��p޼��7M���y��@� ��nT��ӊ^���@\=�_��C�1�x������3yz���_ZQ�p���qI�?#&:4��S�����|�(��n���:) U�r��8�Ӎ��R��T��A��]�{4n�5�b)�*�2�ހ��
���,�\��`pb9�BD�k"��(�ιr�w�9�J�j�ti��*J<��z�}�f��I�C��e���a/*}��)��蚙������!(�iж�n&ȭbz}o3��+�n"E�|"C��s������f�Q����|s�Ô�{ˆ�#܉���`�ڵ���YS��Y=.�p6�ӄQz�l� �"�7�#[����6�t����8��/��+���!}a�1ڄf`a�j���6h�����=]��{&� 2���~��c�D��U<�H���Z=���#K�S��:�-ڿ�~��ϕK�������\���qR+�IZ��Iu�c�����+�{CEd��a��LT�4i
�O����x��-���UIa�c>�
�Ǣ�a�66�V��͐��0�?+
4R6ɒy�ι�@M�����J���>�4$��V�d�{��םzf$}jMP�k8n�
�b��ځ	p@A�a��ʪ-��t\�ٵ��1}����I�[~�_S{��m�j��}�]��p��E�}��TA��gA띣�+3|��/�3���A6��Jٲ�M��I�u��F�A0Aq�uV33��E_�J{�%�94�S�3��+��fLJi�2t�?�v�0~:�L"�,��S��K6��p��U<�	��z5��H��`��Kκ$��c����F�E�:��[#M�.���g�u�f�Z���e)wb՗&���A�u�[��i�\������# ��;"^2d�R�Υ��yR���~�ZK*�K��ǳ��5B�e-�;���b������]v��k'�^��G0��7��R��a<�0�,5Mw������w|r3?��=���D��Q�W��$��yG�^��UX�8*�?�D�t��S��g����#�#���J�������Kt{2��j�+G��*���D�硱R��V9'�N�?�*G�W����^6��ĝ���=���ʢFZ?S�R?��nh#�Ζ��FE ���6��F��B{�D��w ��Ҽ����6&���)�F�=?��_
f6T4x:����1�c��s����W]Ǜ+�������>{�	�i��Ҹ�,R��HN���r[�X|jH蔐M,�]@{$�@$�J�B�vv|������Z���cФ��9�q�J���Q�me�� �W�\_W�����;�R.�������,�c�3�|�s$����I�_�kt~�[2.Z>�_@��2g&��<s��8��}"�&<|u�f��LA��\��Y��&y�3Y���y�ٕ�#�Z�	6��"ܿ�)/	RV7�k�!���w�IF�;��]�����w�9F6���fh�Q��^�LU�L�<9��n���[��=B��HDn0��Џg��qLyܷ�E���V*�����~<YW���K�%~����Ò9��csW:��o�{aI�� �`Ʈ|���"SZ�<��E sF����'cj�7iqGT�ZP�س��!�)/{~h洧�;�� C����vG~,]���nIA`�e$�+y�Z�-����l��o��C,�
7���C�=��{F<������wָ����G��ę�I������Y"~āt�ohU�#�X��#y�N�&�B0F����%]��A�-�y�����V�v�i�:6�D\ Vә��!�o���&8w�v�<�2�tR���Y(����I*VI[�Q�R=�4�W@.���pu*����Յ6,�L.N�v1n)����ѽ��>#�ε��+��o�x��{H��:�	�1ď�B��Pܥ, W:��׾u�4ԍjؑVDr�0�ɹ"T����x]=�:�D���j���j87p<)�2��|Mp*��
|\�+V�[1��.���l񲛋�����z^;�8�p�yXI����zqs��u#������WWp�$���t.�T���ڕ!y�߸i�v�
�r��AL��e[�����|�*�ƾ�Y����Q�-)̌�l���#���b������C9*���7D��̌��ϛ����JG�3�9>�D�Ԕ�jtb�=�<�zSK- 㞥��P%;)��[Y�6�tCk�V}\ ��G�\�q⚋(��ь�ST���k�3����s��.ގ�V5���R�`Z���9�W_�?���">ƕ+�T�yg4�9#�7,��6H��5j�G�M�-�>, -QKS��;�NK����������$�bY�ߙ/X2x�����B�)�Y�^&H�Ʊ��@ ,Z
�,��k+v�R�Ů/�E�V4	���SLK��]V G4�� �����r�K��2�:�E��B�b$���Q)�M�~���U|5��� }�}%X�4�?� �YK�;���G%T0�4e��h��/N��.��H9l���D�'{�Dmr�y?y[�_�i����J�僴n��eg���#���D�$�q��!,�y��(�V������;�˂�K��ϔ��a��V�&�vJ<���Xn�SV[p[�)�c��%�J��{��e���8�w�HE@��ú���j�Os�=P,���+�_n�BBd�˗�{��@Q	ԌZc�Ԑ�M�3����#��y���"�u�/��}�-[�'� �'}$��M
a�㜁�5;}�W��<��ᆺq�Ŀj�p_��j~���(��R�-Yj�Ы)���8�3ǈɈՀ�[�,Q�FI�����`��򆙓:�� �1G���F�ߊĭ��"C'R�^%�������4�j}�y��U��#�P�0�:��K����S�[���F~C"�(	S�����6�K4���Y��d16�S(�M'��QBzw+�ٵG���n6�1̃�d�+����g���� $ڵ3��,ԗ�s���i1m  r.�;2������ڗ�6�P��o`q�j���e�7�m�6�7�,�yHh/��������3�Js�iL���6V߃�YJ-��8-(o*MZ���5�돾�.��S}��k�i�-,ϯ���¿-���kD�ï*�
�Ì'��v�x8�����.�F[�l+fw���/(_�#����z��2ir�m���3��d0�Ҙ��W����߆,��Ns�0I�n�Z׶�~���m=/����w��H�2m]�6'5x�p���А�������h��8�qгN�����B�""���!Ը��`:��u8���XP�N�fv�·eԬ�a��]fh�n��:���#VS�P=w��X�:RƐr!�M6\�O�p��1v0�X�H�a�1N������u��~K)#��I���F���/g=�5�H�>�Kp��9K���苁Cr9����ވ��Hs�h��Hl��lv�ӗǯ���
Q!�?ގ<�eD��E �D~��O@���%gu��7m<P�u��� L���6s8��fqRUҏ���׻ �)���k�P:�V˜Z��ѽ�&D���F�)���F���E=��Bc7���V<(X�M���`���P�VE����c�T�y0ӫ�����`%r�|���$�i�l�=W ��뎍w()JJY��A�z�yp��D���
FFL��2)�U;Gb�ˑ�p `.��0��%����d~�.�\�@�I��O�%�!�ʒ��*&9�%����aY�P�YE���(�'�+��À��@o���5n�Pxs�x0��g6�ra�|z%���}ʠ}q���#鳧P#�{#�������xi�bC��� �$$m��2o70+���3E�Eko��$n�R�a���V�����'%�f��R=��R�o]:ɿ��F�&'�gbQ�RK.��=zLq<�"¡=���'�*�n��n{u2aں�~�Y�꓾�A��'{�܄ef3X�4�W�fF�����!�HɤK[v�!x�aD�����B�+S��Y��w{�b[~���R�tdX�C���hV���Wk+�%16A��3�D�B��#���1��b�3��t�؆~�6�,~M+��0GA�h����)n$���ɨ[
GR�f�`�1 ��s:�U\��k��ڋaԐr�P���@~�4�Ls��<��r�4#cB������Vv��j�H-�G�rT� ���lȹo,ZH3r3�Y���Q����s�}y�4P�m�P���c���D%E��T�G�
�EPOU���1��U�Gl��(?�6MS�5H}Z�{���R��GT�����W���ٰ�Y|~?]l 0���˖�;,߃H�d���=�5���Qz��M��R���
1#���m���jr�}���B=�|���m��3V�K�g%��ߦ�6q���
�5}��O'm`����SZ�)s`KQ���a�Rz��r,��+��*Mr��*HvX���J��y�=`����0���x[�G��G��=���{�����&��k�y�Xu��A�S{�tK�,W���i4n��P�#�b��A�<�O;u��K�KQ���Τ��p��I���>N�yd�\����Ǡ0�P?2�ۧ�\�r�A_�r�dR{s�e"��G�H�/>i�@f9DTdվ`�SI�0.0i{�����Ǣ�P0;]CWZv꺭a?κr���v-h�I7��n�������=�W䦊&���O�z�n��ѽ ��7!�ja��%�ű��v:�*v�=o�ߏ�3��1댂X��?���v!3������+��m�/W�# �B.֌U�v�zqG7���[Z�Z���.�7FQ�A)� �U&���[0ɋ�~��ؠ��\z�v�!}i�rcR9z��6�1EJ�d��x$��@��=�d��"�γ��q�����i�	/CV�AY���˶���c�dx�.�4y�ne�L�JF@,(ވ��պf����%�9D��}�Q����\cOo����ۜ�	�c]��UMB��Cv}���'�j��F/2�$�ʼ5t� �l�$��� 7 �l�S%=����қKv��Qh7g��f�X���4�!����)��t�k �L/}9��k��p�4���b�Dv�؋oM(� �rd����hþS��=T�>��O�8X�ڮ���O��>�0��AG>��z�Zy`���e�QY�}���S�۳%�������7�B�>��L���V�zB?}�?U!B�<�7pbb�wu.����4y��J�Z�hw���� Y�������{f �R��8?;7:��_���\	i�"H�TG���.m7�<T��8I��:-��:P�v8c�y-6U�07sͻ`�'�[�X*/ק�1d� ��������]�슏i�5���r�F��#�H�ě��>G�v��@������!�n�҇�'3��I◙�0?F,��&�[jg�
H����ovx��p����Y�U!#[��2O0̳<�����������D.�5<"#�L����O�]���>=�x��tW$���2|o��K�"l��>H�����GKz�@H�(���@�~�Q��$��}�|j|�xf�I�\�P
]�G��q���2��dN:�xd�v�Հ��ܩ��Iǅ�P�s���ӗ��n��<	����o�9�S���f������������6���	 S-�W�!tS"P������"�x1��:�g�72��>	�m�������#fĽf��G�a��������Xa��c������PH��c�
2�lڣ� KOm�aH����>�3�:I��F�7AK�.����#�7݆����c�鴬@�fv)}���~-�}1*����[�j}�߾@`J�+�,��~:!r���+�Y[���"+��L�nM��#���5�j�uʀ)��ﺩ�r,$�$7�%�)�RF��x����N��3��� <���c�6K��)��_�U�biJ�i��V�Pl��#p����0�������8O�n�-���%(+�e����� "sjj	�kxZ�}Tp\�-¬����Y+�F'*.z����& G� Z���A��"�8#Ye|�'�f����h�8�����'D3����"��L������%fM�H�=Q��˘�|���K���ȡ���#"��*Q���5���4S "d����4!{��T7�m�!��op��D��$�%���S{:{�Ε�<�/K|�pݷ�CYL�-���)o�=5S0F�4ZgJO�Jo�7
�X�U���x��VGO�8��9aá�G2P��7@1����)��1���Ä���*mF�֝�z\#�/z�k �Cx;���/�y��	ǈ`�DCs����s	*����dF�.9Ǯ���:Yҳ[�c�������3��P^T> 4��h, .�I8���I%6�E�+�*Z�e�t�K ��T P��t����Pb�xX�3�D	�X�:x������JR��#�zG��#1|�ppaߥgc�V�~�{���"(� �H�-c��;.V�d���̨vY�4%Q�g�]*o��v��9�q��6.�۩�n�N�u�7�Pv	ܴZ�]���[�����G��X�.A+�6v+��^a�|A�5��;&Oȱ���C�3d�z��{o�0�4�=Q��-��&X�pdå��ǝĩ(�mp�eLk0֌���8��+p��$�j!�l^N'��2�����ګ�����c\��t�CFV
4#lcxN��Qr�g�a���I�f��0��mݚ�GBb�<�ә{�"xF���+b���ɇ�#��YKΨI�s��H쨛S�m�Z��x�P������W��_n���
Y��yk(.ve5�=��eM=�Hý�Ga���F�1P�dKPl�2��e���6�uh�Q��+��J��W?�)��`ް�ʿy٫t7NJM�ұZ����q}���FL���JE�R���Y����eM�VI�	e�R�~�I�M�I0p���T<BGe���t����>L��Nle$:}����@�8�$�{0��S��`9���.�*�:/Ǟ%��0qD!6�P�m��]t�g߂��A*�^�����K�IV�:x�-�/Ļm��+�J�X��x�B��_���K!B*�U�@��b�G���ZI�M.ݽP%�������F;��7��;��6n���V����������y`�y����R@�b��e�j7��ؼfAa��\��	�<@�΋�
�EYz��g5�t����^#南���`�҇�����B�#0=� '�A�ޜ�=4*_)n ��*����ƀ>K������Ŏ'Vx[��@�v� JFȗ+�b�UVUW����[!	ZB����(�js3�鰎���:\�]�NAC�d^�x�����ς�'u^Pz$sb��oڏ��rñ�~<|<]b���;T�,l7��p�!T�E�4fn[{Xx�Ѽ��h�<�#}@y��qm�9"���B�$�양�F�-�c4�l��H�lBf������y�q`vI1!��>X�S�y��;F�ev��U�m|K��s2zu㶳TM�,�'�L�'���s_*"rI�麋~�БtdI���"����K�s �?��U1� ��\������%OP�pR����H��í���'��f'.�ڤM�l����=a�	�<z5����J��N!��po�@:8�L�^[��,�\��Np��"L��~<7�S} ��0�c��(�/t��G�+u�K��s[��d�$��*qXA��ʿ|�Ǣ�ZP߫=X��B=���|΅�������'�0��P��qYs��:�n�o����.+E��RK�Ia�t^��|�Z��@�3���
+��E[�t� �i�tn�%��\I{SiB|M��������5�P�~�3�ǀ��ZP�? ��W�`�Cw�6��~C�Ԇ���!V>�Y�RK6�c�(�0��O��*�K�|�Tz����]�6�ɷ�:�ۼG���96!fR�L��ZX5�J�����ɚPa�Js���W�r�(�7ҥe	���>��3���A��Ec��%� �<Ek�R�)A�Iؠ�p3�X�g�CπO�O�T���ܙ�r�I�/l�J���D������ʼ�➏	h���5A:����<�l�����(��h.���_��b3m��L�Cۉ���U&`NUC�+��G�_)���ĦDSښɟ�;D�]��o
��	B�b⶞Nؼ��_�5@n�w�yDS��	��(���QuD_~x�#�/�{���1k��ǅ���M����U��M{܄�,'�P˩� ��g$����û>P�\E=��!�P��kL���D�[�0�D�ڤ�W�E�&^�{�e�'wMR�T�=^���a|/��������Z�����{pgs�qT�ݎH�U1�q��P����3,�yn{��a)�����k�D�:-��Pp�5��]4�}� t�1�m�ʽ�v�������K��@z����[9T�^��R����B3���A��5�=��	Ȑ����֡y��}�*"�w &�b�{��]�Q$�Ps�!�]���
J.���x/fs.цjZ�Wn� ����/%�q8��,�����#�@S�τ>�D����>X��#N!�Y��4��������j1uy��k��GT��l�'5C�T}��y���mA�I/�#p¤KHA|N ,�g�dKj���5�Y�K�"�CIe���u�H;R���`I+�73�N:@�L��,'i/���!�L���/�<+m��*׆I^`Z��ō��IC�b'2h�TZj�=dS��Oi��3�l���|�
 .-���	e0�=U�hK�\!�S2'I�\8Êt��D.\�a�.�
�@��
�}�������OJ�l�4���	�gf��E^��ܗ�9~�����z�,�"�X���>q,�!W�8<�!��Tk����]4�_�)���ؘSZ������� ���bg��}������_��H��A���g��/�RB�àf	�)��g�!'�i�����|�B5
a[�z_o���6$*�H�{	5^q�Y�~ʤ�cSV�u}��!e �
���z��J�i��	�P�[�d������@� 1P����Xǈ�Y�5�L�Ohj��	8g��\��}��P���3d�EVe�Y���4�k���JdC��\ׂ	�ݗQǙKs*�S�h5��"1�2�����Ն7w��Ų���r���+��3"u���Ϊ�R�榝E7�sM�����?��O%$����Vʰ��ÒW��g��
�	8�C2�O��^�EBj��f�<F�蒐�����zx�mcs��8����L=�z��P�X����V���E��,��� &ͿMfy����M���.�Z���nN}L/�z]-_���SŹEE�����!���Ne�]�=�zZ�Lqca����`$�S]�:��l��5��YkP]��_> �,��#Xi��\DI�0� �⃁���-�I�u;Λ;AF��q�wU֘ R#�!Oݖ�4�I5�A�e�A,���a��ʩl�ע�P٥���O��aW2��ԥ(��s ښ��իC���a�'_Ԭ�< �iZ��EE����)�1O|��n��
�%:�8�B�M�.��	�|�����3!�-Q�x����r�(g�v���3�>`�@�b��r� z6|�L�jLmH��_��3�I���q���*�_]��DKw�a��[���qy͵_S��T�-R'��d����Jn�z�)�9��6�$��l0�!}չ���b�A��'n0q|i$��2|X1�60��x H����p�S<��|^>Tt����o�ܢ����@�Y�#�"�Y�-�vRLӍ7�9���8]����F3c�x$�4ex��@������%J�.��Xc-h�^��r{/h(�0�i��K���7I>�����*S�Q�n��itZ�D&��M� G��ĜD��%��S�$��fk_�8�sF��E��g���!����R9���;���}W�1�K�}���W�O�
Gy��ňz3N���ŒUh'煘p��*�{@=ʹ���y��LV�O2� �o�h�;Md�g����}<�u��Y�0�i4�k�͍Ť��V��.�%�x�i�,��0Q�	�o�Մq���'����������=����?Cԏ������l�����'�xf(i���=a��/J?[�N��AP�J��{+>�f,�CT�&��#*�M}�����:�<=͛<`��ݝп�1�yoo�OD�o
�'�aϺ�T��zh�(�ӂ�]h�k��VlW�ȩ4r��v�X9�>�#t�N��5T�i;��i����a$����}�#<�`ü����Υb���+nUY�ǣn�a�Q�kL@���*���;�0�ߦ�+�Um��TBN��/%���J�ү���o,)Z��W��Pn]i"zM�7�p`��K���CU=<n?�f.��������O�v\�v�1 F�F�Yf����=+�@{oMB��܊H�����Z����J"����W�ڋ	Tp4��*����fy�|Y�E��9�̫4k�b��/LtŤ���,?�_<��ʄx�/g;Nw�I)O�fe7�<����n�𠔺O�R0����L%jpX�U��C�(#�F`��,3u	����sa���-zP����G�`�ڒ96#��̄e����P j��"缒a	�V�W(���*�Ig�s��K��a�����b>�݁���v���ћ�Pkj]r��v�N����;Vr����cic��Ǒ2��yW̗w`�����q2�k�%��ۦ{Ŗw�]�'�D��J��v���^�4E�OI�\\=|Fe��.>ӈ �J��|��H�
�:ڃb�=����Α\?�^����a�J�����dT���l�/�$���ٙ#p�%��t]���Pm%X�Kʮ�_g��P��B2��[�Ę5��-~�()��ҽ�Ǔ����>���!)$><:a�<�U��H�&pz�)��T�Vo`��z?�`ݶ"�-�X9��Wt��ӑ������t��L,N�H�ԅQhɒvu^QɅ�����u�Dj'^�X���k2��ݾ��q3������+�k�I�1�R��;��L�i	agy��*��p�a@8�wQ>e�n���^*�<{ߣ���k!��Nכ���ƥ�:�ai+n5lx����� [aF
�%��$#��F��:�Y[��ڿ�t_����=I0�̉s�ӓq����,��\��<�rtY�z6�����-u���Wu�E:���7�O���zAQ�W�,ym�G�:r# u&�qc��������}7�;A*D��)�BhK�l�^��*�G;k!� ���$Qڱ����P����<*M����&3ߒ�xI\Wj��b�e�p"
~諷�\��y o��{��/1w'$��l�*��j���uȒ��ɖ���)�$u�[�!�RĆb�P�2�=@k!L�1�52HW���L���U� ���|�����>Np�9<-��U�� �V�����dy^���K+��6
RX�9��9���mG�����6 ��s(:�b=
=��]L(�������60}5�q*lJ'p/y�p�����Rj�j���
��/.��[��TK�D�G7b���@rP�}෈œ��wA2�D,��(��Aq7���G(��Fv�V�	��0��bw��.߯��n#42i-�gr�/�@1l{:-b�T�`ub�~����T@�,��ҿςJ�#q���O
�yL	�kD܉P�B{�"�>|p���e?�i�o��w{.z�r��9�7�^<�u1�aF�Y�8��M�i}*��Vҁ�ة5�▌a'�Y��QCiz�{��)~P�ߜ��Ɖ4?xﯸ'�}��a�;ơo�ԓ�S�kٿ�4�8,LD��DN�S�p��?��Qy�S������\R�C����U=D�>������)���sr�Y������P��G�8q D3G��A<Q�/���Z�f)�r}6ʡ/��^Sު�V!��چ��Z���H_�MF3,�'c.�Fؔ�=C���2��ȅ��p�4.�7�l�uTE��G>Y������'�n�Zk���������H��^�EE.=p��<������*;����`���4����8Hy�ՋSG4�=��/��}G�j�L�/�O�f��M[:<}�?)uEY��\x�/_�o?�����8h[gHI��e+8f�[��a�C�*A
�W��绠�,6ڋ�%=����'j��pB�S�z@X���6jJV�6{���ژ]k�<ʥ���YB���D$���:4_�Ǫ�ɵS)�FxK>�����E�����K��ZУ#�!Ҝ�dVO�}�&NI��~�3�'I`�F��H8f9U��/C�>w�S�n�Z�@	�z�=�=�vfA�&��[���.#�S��w{�)z��⚊vkW�U������M�ո����UR؞�`F�k� ,�����<\\Ê��BM�Z Q߾�Oۨ��<�*1�ٙ�Z�)G8�	��?g��L�*Y��v�9COۨ��NRP�UO�߷�䯖�Y��A8,��>C7���R�}Vɓ��o'�h.��+�n r��>�'S���Y�^�ʈF�PW��y�?�����9|� �~~���A'�2�,W|��Z?��AѷS܈u%�q�.e���,*�����
L}���@3��[��7������7��a(W��Ո�?UK��&�=�n��cT��`� �L������ťDK#�!"W���xr���g$�>�;�R�~2m'���5$�w3��O�|�����_���t���(<�� [8�&V�*ZDI�F#J)r��FY{��<�06E:Ɓ�{�<�#�;<�w�%��)V��dU��@ZW��6yF/�*��(�`��Hk����{�V�S����%O�ۻE�����v5rf���SW9��G�e��yâ��m{?L���[״��y�^G�5s�������I"�GtV/�P1(;	��Ni��"��]�|(:j$�O�� ��(��s:̯S�( c�iY��:\h��| |�Xz{A/0����;}V�VĊ�8�d^f���ml��<Ժ�-|,�j����A$�&�b�C[���8�s+o�
�5��Ǩ�a��(���� �pc�xG���s�)�%c�6���@�d�:j�������HX%Q�a* Yp+T�K��2R�;�1(^��!�U	ҽ���}�:'4/����FO��z������'����X]��J���<��"��?�H=�M_̓NJ�5�,r�uIC��`v�"�dUj�$�$z!c{�ɯ���Ɩ�[�܏���L����9��O,�1��7�x��_+�R˳1 ����@ݼJ xAX.6�,�1��G0cp�1=GWr���/e8~����-=��,� ����}uC���A�t��V�--�\i����Rl�HB��E�]Sy�	�m<��������~���3�JXf<D�o@R��J����C:��9>�+�/�IS}n�2�+���߂�xB�o �5>˹�!�]��T$KK�h��+)���˦$(	^w�	*
�9t��H����kZܜ�w5D$��@ʧ��аo!�7�~�%�����0�KU��Ѩ|���鏒��i��v3<V�(.�-�]
4�4�y�R~�XC(��l��_���!1�.W�֎GD?}�ـ����v���iT61�E!0b|�2o`ʖ�l��:qG+�M����C���p��ul�x��tJ�F�g��:�V��2�e��t�2Ψf����<�c��PZK�7SW�XA�����V������U��Ȫ�Q�"]�H1����L��k��
HP��)��YF��� ����zyBӃ�u��J�s͜/Iv���I�6Tv8�+D�9����HY�z9]3�aТ��u@��Ͱ��vm^���R-�.��
1��־"*l�{'���*�}L�D�.+>=�@3	kk��!���Ť�/��^��ʋ��~-͍�v�����v�D3ʸ�<�&��hw*�� e�VcPn��o ?��ם��u���s����cJ
�Ew����F*p�;���x]��u�u!ߞ�u.�+�"�,��qT!r|Q
@7ٓ�,�ԵT�Xh�:��_ψN,s&����\6�����{9P`�?�h���~��mULOꟉmg��׻$��}F8�<�l�/���Ѭ�K^�8��q]@�u��֦#Q�*K������FQ�P'�#��-��p|�WvI�2O[��l�`�])�H陀`�Мyŏ{N����.K~˰/�>=�꓍���U��"�1�ӯz��t�3󊃶�r;l�2�]�w�	���s��T>Lm��@���4����	h�tU�s��v��ϳ��p�~�e�J�Z�~�Q�i#�S�={{�Q��Tf��{/Dr�xU]$"��#%���}������A�9�a1c�d%oN�1�$�R��A�iϟ�fB�t͂�b���#vO}LX�fB�t��7F镽��G�RἯۃB��T=��B�.+*����m�E�s�.ik��-ֆ� ��XMc�LM��q�nõ�5�Q�Օ�}��9	��9�{���"!2.g�/$b��i��|&��6���^;�
kt}F�����l�|i�@��̔ Pp�u�z#�M���ic/�G�)��~�L1��݁^��`���IMxw�I�q�z��j�y��w��ӹ�w��a�Ն��ͬ8}�j��;��p��*c��^u�؅��Sb\ۆ�bƿ�.X�I0�P��oO4��7�W�S�{�M ���޺���K/V\a��quh�jA�痨99�M��7�!�w��X1�k2�';t�]��"�nKm�(�j�a�	�P7#*&��`u���Vɸo�{Pu�%�u�5�<����� �"�J���
+oy~G�����D?|L�$) i���k�BPn#�QQݠk)BuD@�RA�eHF���,�%�����ږ^K_��1���u�'�y�4|B�n1JM��Q��q��wT��f�o]|$��3J����<Q�Z��PLC2�O��n�[
lfiR;�	zw���@E���gy��x��Q>_Tz���Gg^�w?��7i�k�!7�@B����k���5�#T�~�R��&p���<�~f��su�dSa���~N��Ga�� m�'`҉�v�l��JE�QL��@.%~b�I�&�_���v5�d8���v�є�jKb0B�Z�;��Z�ME IT��ywP�U�W|r!a�"ƣKl��7�LHF;m�U�e}�$�{��/�f��1Kq�z�M7e�8r�nL�8R�йc��}��q��d�?�U2��9ۼ���o�i��U��ܨP��4S�x��C���㽸m�^P�|q@�`v9��dj�?�٣4�0��^ڜ[g��3�h������/��Iq��L2"��U��(��g뇳�_0���4�~��i����?�8�?�q�u�t^�������I���F��߅&�N=s��Ԯ���?*@1�N@��	��-2���oc�&$�y#�����-�h��!��flK"窜A��f��"Y��l5aLy��/�=gyM��%���S�>�4��J�x��r�'�ds��?����L)�==ŀS��KI�G����Ą&f�7%-��bpp�9���dʑ�+��K��GY|8��	#�r(_�"�7��������'xջٱ�� ���+����q���4)k��C�8��l�B�ރ;"⣂:�|J�[T���h3����S�/���jz6�ï����x����9�����X�}_��D6���ڞ�t9���t�=m[���oH@�S�%��FY5�T0,��戙͍n�ݑ��%�#j�� j�d���_r���*�;���+$��9���E�fw|�ý)�m��v	9-����i33QO�-2v Juк��>O���^la�?(pVs�/r���;�� ��g}#�PrHu��m5)��%����L��#�酶�����\���,���A$(=���Sh��V��)���W�[]�T�I�8r�P\�9D�ۧ�ֹbChaG���O#7�rD$ߐQ��J��P�L�Y�Z<�jx[�(�Ϫ!G���V^�4�����g��C+X\�J���x�o����3	u��7�B�E�Ö��l|�?�UF�ъ_.�t\��`�ÑZO4:�:X���I0�!X�� Q��QJ�P�"�漊�BV��`Ed0�H��)�Wa�8�L��Isu����1�7���L��ǩIRAy�P�&�mT����`%�=��Sk���?���F��iS�H�� $��:G똔\�d�fw�D7����@ N��}���㗽 pm�E�ªm���A{����X�0*�| _�[��� |.[���N�ol��Sr�Iꂗ��0�^D�U^�TD�Ӌ�7�&���"mu�\�͕���rQ���Q�����O�K�%T\D���"��c���F������Pa��S@&����X�B�ql�J�\c��WV����oXڔ�����tq����'����b���� �o�y�p��.�S4��ew��L�t�	��#ѓ)���9�{ ����y�xH]�Ƽ�<_h�~u6J��RC���.�¡f4 �t#q�a(85fIh�	�0����b��|�n��Q�>��T;�NS`�w�^�/�l���A����|�L-���)Y�ĉ��U�@�#\	.G{k�G�-�;P��͡sj��N�#0�!���ψ$�EDz�ن�\A����T����K���&��ԼPH�o���jw�>��;x�^�G+�P����Z��U�!�B�;���t�B�ֳ��Q��h�����yF6����쳤��paf�b���9�!�Ǎf	���x��uZ0B̟q�&#}>�*�����Th��`K��U��!E2�W�#�+=��*]���F�[�#I�fیÎ�e����r[k$��ban7l���4�6*�%Y�IA��L�SF�#9d4�S�Բ~'A��%j#��$�
����o���<YE�yϱ�@�D���L}Y\DW����*Dvձ��MZ>��@��g]�YS���l�"�$�^aCae�+A���l���'.Ҭ�+�aT����|Qe+���t�{Mޭ)��ح��	���_͡��ꓥ���'u��2�eH6&�C��OBi�;s��)q�Z� �z�).�8�H�>��7�4�O��t��]��{
/����Wj~P{�6U5�[G�0V୩��]�{B'6g�\ Ӯ���6���kD��i#I>ZӜ�������]jw���<Пf	�L=�#|]�i<y�������\W6���&h?��04�x�D��4x�|A�sp�q�\F��lIU�����]l��mΣ ��Y����p.Ϳ��	R2�Pb{N�H�Ri�������K���z��c���^�W�/]?(���+B��l�8�6��#|��V�z7�Ig�4��z�#���; � �,{�8bO�u����'�?eb�I�[���܃E���da56��H�
�I��R;ix|O��>h�<�T8#��X�>3?à�^���S����H�-�^�V:��H	v��kH<\��H�ͅ�Mm�R� ދ���.��xp��]�)Yp@�l:���>��t�{# :czsr�봤׻�6%�	k��n��HX� дVG���b�l��Dmd�!�J_% W��q�&����ȃg�x#�.��o'묓:�h��m(~����
M~G�ޓ)ZVD����N�S��-�_4m*T��s��g۶��F+��H¯�(�x/Ԫ���&�]j=���~����߮�q4$�$����B�z%�����@I��k%�mϦo�`����%ˉ(��(H᲋�\({�c��`��2PZ��9����/��͞���!�7���TT�O�H���B�o�@ŋ|~�eY��&�u"�N52�7�Љ%Rn�->�� �J�W���)�Q��3�}Cokڨ�D+�X��v��j��S��*�*I�)t�ap2��.�F{�h2eU�J?��>:]�$�-w[Ms;�B�.�T��������i\�E�R~��7�t3_(��΁�#ҵ	�^�۝9_>�T+GEk�$g����z ˎJ(�h���{��i���?#�ޞ�}n����r"��|;	Z�t��3��[��7r[煾	�o��J�����G���t>9`bsP{��<��}0����{;�ԛE��$��F^ui��h\AV9�o�����z��܄�f/�8�>��5f{z؊���Y 핛Jű<>� E׏hǽ�g���ZY
j�XϨ�2S�T� -�!�O��2R����b���ɮ��3əS�x>!X�L���]O��h.{��g��M��-�}/�ř��O��_�p�����́���t)m�:���8�MF��x_���M�^�	�@��y�aV���7H�;�{�,����ۈЗ0n��Z'}}� >��"L��`�3��8��R��O��2PjX��Ć�^����-5��v�L��)�W���Z��deQ��9�$J��@��z�s��c���%ʽ"�i�>Us9��%��[|�hMF���$��	b`�W�:r���qg�7��_i�X��2F���"ā��Ii�q�&��ŧ���_�RKN�꡿��U᷏S뾤]���pI���6y҅�Z�_��T��$� ��Z�����*C�b�q7P���`�="L�X��Z�!K8�Y���R����<6��iEI�lg���4�V�>"5 ��Ir�1�$o�F��NW�;ƃ����+����r�׃#Ĥ]���%����L6&����9���!�ڎj^�LI���fwԢ����8�*}���Z�/�P������X��n̈
]��O� f(��-��j\橒��-`ƀ����I��Q04h������[�\���C�3���,���v|��W�Ge/���!0�K4����6��U�>��tꉉl&��Ζ��k�H�0�;�I����b֤�g�����i2E���y�D�Q��]�_�(�t�E����>�Ք��U��)�h��^/�c����)a��U��.m���zX<�?%fF%�t%�D���/�6-��´q%��a8�p5�A�gNr)B�|�ȅ.=�"OȻq3�K�0%��T���1�Fg�;kJХC��4\�'�`EG�LNX�4u���-��4��c���`������zl���Ґs=��ZUxf�g`k1��}�"y4���q|c��r�|$�����n�n'���b��.����
��b
}�S��0��o�nی�͝�oT祊��J������{ ��=�{x �X���	Tʆ�p�wJmp\��m��,��ry�\��2pW���(%�ᢷ0B�Q�{�����P}�D�}��(e��h����a;n���;����{���Ḱ{D�X�O4n�<c�
ۮ�p��#M��H@�΀�+�zb�o޲�u��M�u���(f�o��m^�!�dD�-f����	�&|�6n'�U��0鞆�W/����W__z�	��+ �^��zc�~\�X�4�����(Æ��8#��}[�HP`�T���rJ�e6|J �j~���Z]W�S�����!>9��1�D�J7(�gi�3��`�;v9t� ���hݙS�y�)�����?��8���H�C����cJ����-���m/� ��H��4}(���c�h1I��u7M�[���D�ږw�`V�Ќ�-�����s�Ёa�v����/���~��3"݄���}w�-x�=%te>x���C�P�?t���d>:>9�eCj�+Ttצh��N͝Bl����3n-�+��;c�%-�Ph�N��D�B8�Mo �6�(\ʬfS�[i������ug�GE�my�~Ciք_��= %U���BR�9��GK����<6Y�
1ᣛi%�:K�+,:
O�FS��,�EX�^kwܪ��]�F��#xkH��.���c%pÈST�*C��@�Asz��K��<f����L���$�@��h-�d<�=/����	K��ǿҊbCx/�ܽ�5�v�R^�rr+IKX���6��{R�k�4dB]u�5�FX+ �u L1^ϓ����h��JUXOmJ�1Ӫh�]���e�_�����z��B�L�'��T'ʾ�-|l�o�6��¯�/�`�pV��	�о�ܘ�����"9�m����z#�³�����9u����;�
��:>Q��Y�ms�Vn�E+�!�e"��n���ϥ��1PA�s6�8��T�Z� ##�fʏ��D�r�IV���3�w�*��R�(�0@S��&��fsl��w
'%�>���.������ ;��-+�p@�\p mE�2�GXeta���^B`&�	\r�|�`��o�ty �O �W��IP�������fYl�u����Ch��C$���Z<3Kl���ߦ	��k0����H
o��b��@H�|�Ӥ�5�X6��������5l�G.^���vMa�K�y3�N�X��V��v�ߧ�fޔ�'l��3/��[���^!���t&�������� ��pL��fV;�s8�ImCR�b�4��.�;r\Vhq2����s�3$�E��p1�Ei7��'G4�$����XZ6DM�Gx�|PP��Peʔվ2���7�2 �;_��ͩ"����4%�D��F�S�כ%�4L�	�q>xޔ<@ۧ/X�x����(sr\��RNf��5��n��8�����y!����G�,�tn��kUت2��b���`M!1x��SR��pq�%���s��k��*
�����&�u�좣)ȶ�E�]qP<��^
p��U:xvH.�y9VҘ��Pp+��]�����ν{�y�n�1��z8�,2�0FB�T����<�!V�.���V��͢!����|����z�	ϫ�ڿ��a9�D�t��ma�L}m>:E�0#�yu0Y���p�{r�%��2 �'	`-��}4�/��ކ��)��Zu/w�q�I����c�4�͸O� ��|(FfW���۳��p':��[TV�Z��0�\+��)ILT)�C�1��5�G��(��O�����r��	��Ahv��u�x �����O��*�8E�L{�����['�7ϵ-u [��0MZ�����ź�t5.�3��Ǵ�J��M�6j��1�����ܘNh��>���JW-��d�:�
l>�.4bs���#Vj�г��奔>�͠�P_�l'�,�.���z�Uj��޻A�ꕢ06����2�gW�9b�ڱ�foO���kҨO��dj�������J��!�b�ԍ�*[�|����J�^ЍD����g��\�WFFsc�Z�
)e��JE�$8u��w�		��;OZWp̘ra����i���}C�^+gӂ����ǖ�^Xʏ��N�� ��X���М�[�j�������Vs++�w}+��ML����-[cT<�g:L>=�%�}���ڏ��Z:%,�Y=O������1��r��M,��I'���l��f��4�f39��΁.�Zs��0�
|b�s�w������:�g�W�_�!t������̑,��A����`�^�`ev��)L��!��o������Z����9�N�@<���ʞଷ��P��Y�� �kc��������'��JL����W��M����܎�z���[���e��5�Pv���� ��gj�0���{�K�B��',�%����kd���3�z'�.F��f�[���_�����v<�t
�t_j�����rq�~�7e[�Wp/n%�y�����g�Ѓ"M`�����L��ldЏ�ٛz�Q���@� S.�d�{.:)و�9��"D���qHQ�q��:R[�e\�uH-��bS���p���ޗ5���y��n#j<Q����/���]���a9>]k�-}��z��V*!˨ͧ'�x��DI�~}l�fɋ>TJ�h[���H��?��r�=\@ې�zU�	r��XL/������#�`�2��M���O�M��l�Q���������2�F-��*�mo�����ݴ�Ru�W�t�o7q�ǲ����NK�<W֩R��Gٞ��_���<v�	V�#����2h�%��\WD�G��"PIo֡��6h��
����wɎ4Z���٣�T��A���PL.@11�e��+�0��{Ȟ�S0�������=�H��.�k���8{'�m�o1��������M�8�ß&N��f�D�~��!I�����O[���U'��a>F��'��
�ۣP3v��3οY�0��S��l\~�g\>ߏ�źׯ�	.�`[��v+�1�*�Ph[M���֩l��zm��#SVH�(,��E�1B!V�4\]�ݠ!��z /$��@h�rl�n�?]�Z��>M� I�P��@�?r]HMZ�7�7�_U��t�j�G��S���ƅ�ߙ�����p���#��;q�	z|	����75J�ut��)���6��*��*�
޸R�R듚�0z�3,d���0�C�����*K?)_��h橉��h���Ge���^.?Y5����
������}u�7$���¾c�l紊���}s<F�����JZ��
���=@H��i�������G���+�BH"���܅@��|0�MP:�����p��6ob�;!���G�yY���QQֿ1�v�/m��|K*ý�����?Bn�`���|K���CL[�����AG������&X?DZ-h��r7��� ��.`B#�	b���_��������u�O���@�JL��iz��nSFR󯄳m�1sx�nk�N�`Z�{ �iNw����f�f�]<�r�V�~[lm��#��ʱ���m�E/{����	mZ�¯`s�,��RC���g��\���F��f��[Aܜ�l7����
q��)C��h�t=������Q��n�4�s���D��k�}�%p���,�6:p�����drt֮��i�k��]2 ������8�K�����Q\
aԧ/�9ݽ��5�8-������۩=�[�O:��=]�9v� wN�r~���j_W�����0�!�c��9,� Q������Z��\H
�?'@k3�o#�A
4]�C�C�q�A�,X���0)��Ɏ�.of멃���?`�b)/-������SC �ȼQѩy~Կ�+��[;tg�u���!�(�2�lo�D���,p���d?!	�o�_ڔ%A�����ҿ<'�H������|�k'�C-8%N0p�����J$o!tG�?Tc��ݐ�
�@��;�"p>��Ň\�F0z:�.	s��`~�&��˔��+���b����$�	���_�]��L�>|���X���~4!����	��ϭ-�4�q��B�E�SHL�j���&�8��8VRK��tNӮQi�|��=���3V��C���(��}V�bQ�<�-g���N3vA�Ȱ�#끃P��Y��_�� K�j-kT��^���|���$�h0x�Zk/8�� D���:�� \A�dnX�G'����ݞg]�my�-��GjD1)���#h�tYn�$���6�y�'�5nl�$[��Jj�!���J�EU�ϪLu���R�!�F��>��վw����q�5e��_�Q��2.��)ߨkx��z���H�s��i@H��Z[	z������0y9�j���G�8),��c>�xӕ,p<}���vz���J�$XwXB���V悥%v�Ep�t9���s�Wyd�.y����;�\��M��j��.�{#J;�>:ⰎR����qM�(r^R��pK��Zoꕋ!���!����zX�#��4�&mD��!�#N�W����<e�{.�2U�[���A`�e�4)�XK!����z�L�\��%�I�A)���!d�R�\́8����Id�{%�#+�=��ɠ�1`��8�&����\��A�[T/4:�?k;��z�R8�3���MO*|��UG�u�S,T]�.y���7ӽB6�%O9Ť�����z��sc���u�#}���Ƿ��a���$!�.x�\&���W�QJ@Iy�)L^�!���L�X�u�?�sa����}�-sk1��"�µX9tv�,�H"�$ `�u���Y5m���˭
����F׷6j��"�*�~��Y)�6͟.?�"�Gy�mf]��s�I!��0�# B\>����/��;Ԭ�˯�";��8W��4���(���/�5�X̔ݪS��[)d4���6�@7�qh'J����tT׳�a��E Ս��7G c-��Z^@Z��83�Y��=��x�I�Ч*�EBD��p�v���ԣ���Ĉ����46�K��&˞|LBV�W+�^��t�mv��(@a�طb���p[c�r����+^�PmDo6���:TD*�A6f��?C��ۉ	��\r�e�����-�r=��#m��	X����6�����_@�$Y���4�����)�0W�kM�_���bu5W�n`$|ѓ���� ю�"��LG�� IF2v�J�E�Yh{����_�F����g���q�<E4�o�J]1�`]�_a_%������ٝu�4U�HY�M��7�0�(�OѦaE�>���Y�Gƛ�u&F?��j@T@�J$��Ns��E7��=IFl������ݩ��)����Y#�;�;��e��VE�=�V�(�]]�_z�\�a׺�`�Jw��%˷^�7�9(O=y�h�����P���{����d�l;�	cПr~��n��",,�h�u4.����u*�D��eh�j�|H��7����FS	M�b�3"��:��X�l�k̢4��N(��.[�5����!�{��wf�+�WL�	�^MnmZc"M{d/[D�N�64䌗Q��w���)��x���H�%�N���Ղ�{2y�!v`!��\	v��S�1�����o���0��m/�H�}��P|H[������B��p � �6�"�C�J��t���V����X�V��"��)y��~W�*ojHB?Ӿq�f���_&��h�eŎ��x�G<C��Ҩ��C�K,[�}��U4��;����[�����1.��i|���F�t�s��Q}&a�*SP�n������)1��qx�ӻڸ��������OE.|��}
���� F�pC���y맀��S[4�Y�
��]d�e��8�?R�?�е�`NR���� �&�i<�Z3�o�[�n�\��5�.��ђ
<v�k�	X��L1�5�Y��a,!bw��k�#'��@���,c,��X�f�[��֎�}��oZ#�^Xof��b(�.��N�r,G���X��6(��|P���#����İ�������E�8���U򥵾e:�9�Ի��Ɯ��m�e�O@��ۼ�?.o�z����$��{�B��
�W	{�|�vc7v9�M�@���w˵I�m���e�x�8Ci�_�X����0���:����sz0���X��-����i�k����*��)����7*<W��r�ds�Jȓ� w��n�)�;����\H	 �����NY���� m�j��KD�&�e�-�����-��72	��� ���0m̒��0��פfm��Y���i��9��=}^�u�'Ӣ����@G�x]e���������ag��<j	zn�rWgw�����z�t� �c�q�n�:m�l<~ƽ߅B(a�[�Ƨ�6�1�q����"`�Y���1nE=�����#��ۚB��X��~����a(����9�J8;�L��ݲ��0�<��)u�Ɍ�����;�·�??�Y��i��S��-��N���G�A��<~ йG��ʌ�+� دԞ��S�,zd�#�ŝK�H�S��K%�F�W!��x�!Υ�y����H�5u����~k��e)�DC
l��|��n�Gg};�3�_"�1�c��4r�d{���A5��!��]��i�Byؓ_�S751�H�<�{ܥҤ�c��{h��4��w�����R8���~�8�Yڭ�TB�x�3�=�Fށ �?�̊���p�gga1��X��W�a}���e)�i~[���?k*�|��q�
�zWR�_��7�D[�^#��.���@h`���ӯ�� �V6�_Ȍ�EO�?j�FGo�������Fur�))n��kr������}d���K~�g���(�*�8z�����k#�G��]�oF��j�9��`?W��9�Qڿ?�
o�,t�3���b�a�4&��9���Y�'���������*i���]Lz�!�f-q�I)|��|�hI�5�tfh�k��_�%y¿]~r��#���ӿ�ǉ�-r���&O֪�]���m��D|N"�&��*����V'/vJ�h���,�ٕ�m�-�ٜ厑B9:���n��ٽ��I�H(���A�J������h�g�PCH3���3%uё��
�e���v������!ə�-������@2�IW����}Z���y�ϛB���/�����*��0N�*���z7,P/����+�D�gP���lO4t�a��>A���|��!�cŤ�o�l
^^R3�9�ƀ16gyƘjϣWg�����ӱS�p3�x\�sL#�!�&�D�}��I�"�?���Z�k� �o�eNp]�n�S�c��fb��qN��B����Vթ~3.��{��r��*1��h�/?�
���oȤ�I��ɷM���1��Ҁ��~�4|S�Ѽ�g��#���#jv��>M�$��w=��aN6?$�(l z`�%�_2Bz�����o��̖yp;�U]��Uu"��J��ZsU�"�o��,f|�h�� ٖ��	S���4nW�hRy�]����Q�
6ń�Ѱ�iЮ�l��4J� �d����V�5@��-ʻNƽ�~>�(�%O.%�ի��v����%'��!pS��Z�0ρ��R��Z��X�i O�k��8�J��D^��J1�ZB��j͓C��$�?s��*c�f%�h�^'q�9�2�5�p���yh���i�>��9+ݥ-��R��+���/�m�R����_bۘ!�%�O�L15�ʥt:E��"i�f�u�z)���#=aά�y��2�j&��?�N	h�+�� ��z�S�P�4���~�f��4_H�4��^(yK§��1�o�a���T�!nޘ�0�OxL�jl?�d���ic�!��~)�nc@�$�s���X���3�L��C��L�m����v�pu���4K�����#*յ5�%�V-�[?����y� �c�{=i3���.S����]73�����?�j�k���V�C"XVN6�U#b���B��S�{�1���V����)�n� t�3������/:x�N�`��Kz�M��|�I�Yq&u�!�,����y���g���1�Z��߉�T�Ƽ�*��`d7$u�&��N�0�ܲҜ�X!��M �YfE���p���m�h1Ƥ٭5T���oDd5��c�T�.�M��}L���v�4�$}ӵ��y�l����%S� ���@~�%]"~CIc� M���%)�gs�u�v���D�WP6��H?�@���i�;&�Wh�����]b��y[m$��̸)������m�g����-&�i^k����V����S�� (6sUr��$�L/�]!�f�F�C�1@����R}�^Z+ڬ3�P���Hr�;N�t`������8���fn�W�O֞]��~�.`0�LR@(��f��όG�[Vh��c� �%|�e��.1��T��6�@��=�5@|��Mh7�܇Q8`�
ΜO��o�|�� 
�p��۷���@V�Ux`8lU�j���.$��|9t�^� UX�5EA���M�|S�HPc+���y���s��������@|SfU��Q�/��p��B��؃�9#ONgQ��4�K�?�eO0�����G�:��Q�N�#�e��#ہ�pU���%���0ǸgO!7�l�\�m�({���C[�T���n�0��i�e2G/kk���K����9���z�:��9�s,
<�Q�2kƴ�{�k�\E���%\O{K�7;z��j-{��]�_�W{}%�H/��Y�V��!���]�5�M��>h�\1�Л�O��4�$�S�f�ۚ͋�RC;\��]ōE��e_�p�8I��h��΀/�@Y��+)�պ�%��R�q"�Ke=	����^�"2h��ɂ6�X^d�����¶�1{��b蜗P�� �!m+{�D�J3sr�Ø>62�SG����׋� �4h�8Gu�����8�y��d�!�K�hP��V�@K�T�\��N�{�NJ ~��>�3��#J�Tݬm�=^���o3�Ѹ|��������$�����K_��ّ��~UU���!��&�N��z�'�E�Z蕬��;�D�n��T�yw������������q �'�����Ǵ�1C��L�ޚ��"qɉ�Ŭ�2m'�Uȓ����xg�Z�'�HA�y��w�����њ����������jQ4��a�
9V\���F�~q�sl�9��j_s`%O.:U���lsS�n�.9���R�|�phV�h�J4����s
c�`;�R��Hb���z���-w2��D����]od�8�HΨ%A��L��W˥($,*��QB�l�YCb�xaTC�z�	�1�s��2���[�e�ܬ(M����A�Z[�QΠ���O�M���Cm@�<�%��F�){������Q7T0mõ"�p���O.Y���J�6 �{�!S���2�6OFO�/@�2��&�Rh�u=�� �Xh���^�I=Z�O>�yW�V�q"�~�s {�O�5>�&LY��[���ڢ.%�2���VV��3��[Ƶn��P$r�[�Jdw�5�'y�>����{�^��?c�!r��6��V�d���86�`7v��du?
s�q�9s����㤕��5	��'�~�#��e) ����hB$荾��S� ��c��o�:9�ܵ��\{�~��)�\���@�n��n��Ů4�c�4C��M0$W��ݑ5�V�]B����<qD�C�O�Soa����z�[������0��5p}�Y�Q�^���{H �qT�&��ʦ�+�7������V�aX8�ԉq�EKý�N��Y�T�Ϊ6��L~�0�\ąAg�g�8^��<��_��_�A,��4NO���g(��� �.����%`z΁��C=xl�;�����=6K�7�hH��:�t�n����<���;�������؅k�=�y��ϯ=��9�+�*�P}��N�A��75���k0���慭��B"�LO �4�Aa%}F~j���U��s���*+�g2�|�[N_�F�(.6eSW{�?:��V;� T������7�7'��hY8������UN�h��`ے��
d=���1�IfDY�$2,&��'���O�ҚI�wz�кM�am�)��&���B���*�o��%B�}����~g�(�!�Z@t�1���՟��Y��/vَ,Lޮ�JzHId���"a�ܗ���$��v.���K��\�<ޮJ��wms3Ŗs��u�+h�B��l����T��xA�^l(c�3З��&�@�j�[8~�t�ۤ?.�m�h��X�ֱ���� ͯOپ@�dXq&����)g6�Q�r!����P�ע�]�����b�%�[E-L���Z�pG�����KDLy�䭧j��OCM��P@���,f���l��[6BW�2��KC��+.�"�P"��ԫčq��b��*=��U�{�@	���˹��qZlM3���Ρw�CfL%��z�,�nY�כZ=F�5�1�p��Ɗ.�Y�>k��E(����p��R��r{/10�I��R��ޔ�2-��H�\��qr3�ZT�&=��N�晪�0^�����A ��J`U�E0�#�[=?!L���"I�/0#�RȄ�CY���u��������a�G��HQ���Nb+� /�X���NvhO����������KL���}	C�r�]ܖ�n�^���b�$�ѺI�1�o���5��jt����1��,�	��T���_t� �I^�1�ƫ0�{.d�q��,�q�99t�l��5�q�!�pxNm���3]hu�.���
)G�%55�����Ue�U�Y�K��A�@��5�e>TdQ�b��vT��rM4Y���y斉q��>�0)Pl�v8/�a+��<�a�v5�_�V�jH$l�|Zy}c�X���?}��@u���5Mc��DM6Qs>Կ|�� %�}�}�4�5'�^C�A��w�3�W��G}5[��Dn��u�=e�k��?A!�څ�.�*��g=F��?O#��W`@L�h�j��ɵ#�!�N�%�.o8�pr����>53$��5]�^��*�w���8EChW�lJ�D�� �9UP��Ɗ��0���X����� �K��4�]�o�!Wf������/�S�	!��[<���4f)3�Є��3d�x�)ݿU�v��[��<�A��n��h#hr�8�
h���.�wA��8�̭Z4��E�k^�)��G]6('l�y$���כj�|GT��T(Uw3�����p�E8�Ȯ�ڃ�s/ `J��V</ʔ�`-��@l���.�$r�p�~v���G��o8|�=mѕ9G}�`ֹ��e�$W�Yy2�F�x�ۆᑷG���@�Mڦ"��K)מ񹄧��;���M�S�����Y	b�*!Ht��v��w�Wzq�*7y�1-�դ���D� �r�'=q��������v()����?C#���� ��PZ���������m�\�f�Em��Ԁ��{̏2g��I� }>9�S=�8��wU�>�e�#S˄B1�N׵��~��`��k��b���G>Л�\6��fU���h�S�Λ�N#h����mTx�"b�b�{�,���\���ͧD��u^����TI�&�6��4��5����u�~�:ן��m�������q�~�<�K��]��(��Y�kG]௧���ja�b����f�QE
�R@t�׾�n��'�E�2��s�CL��"�Q�����G�J�W�{*�E9���Je�#d�%���J��3U�V��4 ���v��Dη^i��9��S����(D��^��ڄp��U1&��ű�����e����Q�L6^�M��I���!� �4R_8�o�K��O�_��ǘ�B�P���"���q2�߬tP$����N�Y+)�t����L�,?ݝ*^��m�m%�Ў�Ɵ��*��h��M;1�4�y����"�J��[��EAS�wǱ�7a��7~3.|����2��xI+k��1X}/�J�<e�0N�oRc�;)nD/vc!lY����n+�����OpJ)�4∜�r���v�R�@���O��JfGL?����Z��� K����+��k��V6����M���g�j���1��^$��)]Ѵ��f��qҝ(��5�oB<�L��WV�&���т��m_�1W�e<���,�i�^���!��c4|��A^���y��n�\2Ch���9�[_ѥC����{�yu ҝ�������佱c�����f��p��j]���a��\��O:IS5'����]o;虸#��.<koL��I�&o��̢5םV0�]�b�aD�H��7�M]c���ń��3_n*y�Yʘ�Չ ����L-CQ��$B<�>uV���}T�2*��9~w��S����DG�hř��X�RbsN�m���i����ݘ7-�Ѐ�;��qNW~�k����s.tĨҴ��Gk�4.krc�z)!��/@��Ѕ��`�NS��چv%<Pg�Y����?�1k��T�W/�7.y��P�+i4�F��Dk��p+�Q�j��] �����������i�Ӗ����t@��M��92��R(@�00zH���< �����պ�Az n�4#Y'R���%ɑ[�)ձr����,>�؊͘����m��K{	��{�[���1�Yf����zP����zٴ/n��TZ��6Q���ʫ�F�����pY_���8Z�,�pZ=��C�� ا��~vȰ��@b�ү�fJ�����1�{�$�b)���j��e������@p�Nڽ&F��Wٸ�$ܫ�1a����c�ϤȀN�r���F\�&�멝|m��@���)~����YU]s������`)�@.�?f��O&�~}�]�5�_����Rݚ�\�T�`��y���:��j{R4b1�����s�(׊ʡ"l�3�S(���{Tx>�x
�_j�3H���=^u���M�T���2;ؚ��� �X��o���>L.͠�QO�����?d����=G��.J�i��>_(�K��+m����P�'��1۽R�Q6���R�0Jo[~����tj��k�Z��NX�(Oz���C��B��3�G����2���� ͓UH�;?���x�S��qc����ND{�	F� ���&��;��4�����l���j�2+�� SF���xl�2��
���N ��8����N�A�\)x��%e)BE��D;��rfO����M-��p�8������Щ_cٚW��j
h����=�>Zyש�j�fE{'I42uq�"��Ss�4vx�Q�z����Օꂇ.$��2�����7P�l��5��2�=�I� <�<��2���=�I"h߰U�� �?�*젦�����Q�\�����A��ԥ�m�Zʣ�G�o�eHm��9y��Ua�=�Sڎfhja��j���j����x�SW�2c�KS��W,92��I9�x���FF+('�6��/@�A \)�"$ٞ X�*}� OB�D���KL��a�5/k�o?���T7F %��{@Q�;��M�����|]�9_��<~O�0�,�r??����h9�����rG��������=J�e\����c�&y��a�7g7ORo��sŽ���P�ՐB���"v�ϬBo���D�J<������;����л�C:u�e��i���"��jH�O��aK���~�%��
����!��(��1�ȽBM^z��O,�
��i�N��(�_v�����2K��K:&� ��RQW��>b��(`0��z"Rf��NPe���5����Z�H5��b^������г��S�Wi�	�Q�h�'�xJд8����[�]����*d���)v����4i������_Qh�{r�v1d�9� �%�Z%���u)�,��ؑx{�.W�6

�i�B��u�(�u ���0�P�WW� �m(�Ѩ�f�:�
T�"D�\W+sL|(5�K�V�f�拓m����)��)頟-q;�X���]3�����+��Q�z��Ե��<ĥn��%اB2���3J�#���w��Y�=��J����`E	� [��a�|�N&����GG�d�1��g�9c�K����q��a$Q�	v�6�¤���&=�R�]�܎]х�<p�#�k%�L�摸Y;1$q���ϧ4\(e�H��S�J�HB�	����ʀ�;���X����5��i���M��u�O��Aw8l�$M��z� W��\�~Zs� �=�tN���s=o�֕�N�g�͐�9���8��p��5��f2�B���>��_�c�@C�QE�q$�~y��<�;�Ci\5VV�0�y��xYbv��4
��t�M8O�v����-ok6�75R%�5bc��h����{�#�CQ��H5se�੡����3���UO[E�Z\@���*�ϝ:
1�����`
�Qa�}_Ү�/{,����щ8Y�w�Ma�Ah��Z�N�j���5G�)X�$���@���6]�3j��� 2�Ŏ�gI�"���mQC��rޢ�MmX�R�c�� >z��IX��sJ�x
~ ]��=t�(>X��^�o�*�J���vYC�@�N�mw��bU�2��͉YH����V�aB��o�EI�C:O��m&��c10)�H2ҋ!�/a�����v�Gg!��ٙ#�1��.)�^Kg-e���!�'��[)�Y܈�jlC]��'W����ND=����k�$ �%Hr &��}�rv�b}��W�,N�Z��?l!M��`�{<*�{x����,��h-�� 2����a� M����O�v�#�CƎɎ�OZy�MX�Q�y�9�G+������^�W	ʟ�d`���G��ĴQ�x<�	" ��E�B��t����͏�==H��ƕ �䘞�%O�I��?.y\V���z�2�+��Lʗ�P}�����=0��jwV��ˌ�����O�mm����aPov�j+���\U�C���oN]�4|�<Y�0��~��b!�W���Oѿ# �'�s���w�Ɠ�A\;��E>�w�~ �:y�)��=�S�Z" �%[��+q��G��oEZ��!�I����B���[?1�]��d��<-z���XȤ(l2�y����V .�C��2�G���:��K��D���7{z�ƿ$�"��\C�5�fp�c���1
���5�e/@�VC}JD��UR?6�J��C0�iX��b�Pw�/{r��c�H����Z��z�@TH3�X��"jԓ�X�eX�Z�n�������Y�0��������z��={;zR�|s~p�����Y�Q��}�}��5�1����f�p?��
������f� �.�*��� �-� \�~8��_�ʃ(�)�O&T��a`�?��T�_9K���P�灨�XT���^�����հܾ�`y^xH��6��l{�͑2c:��ʄ�ƲY�O$(���j �
��5���Uis�N+r�w� _��ڞ�1��$���g�fT5�wmS��ǚ�5\~�;�q�[�?d1�0��r�82S�撃��$
.K.� �TV0�p"���m\r�.�*bb�Ϙ%.�6��h�x咻/$��Cٔ�e��ӥ�����Vkʍ�g�wV-Q��E:��l��h�` �&��S�#�z%J�F��>��4T�UA��oF߂Tq��W����@�E5��!�{<g�`Q�
�����o��Z<�
��^՘$���?6_��8⟛���=I����2H���5I��x���m������A��{_�����F������պ_��7uù�7>�?�::n��~5<�"k�`�$�j`:����4����ި�!ݷ�����"~wBY/�u܎l�����۹�N����L���	?���1����X=w&��5"d��J)��/_ T��Q�|z��{ ����`L���aհr��>�H�&�@��<M����Nt�;幈����I�V���� =R����ߕ�z�>�ϺJ�׽��^q%@\o��Y��sb��n%
���&a�G��kEz`������lwVI㻬ݲ�<E��(�Ul�NRQ��IDO�xm�8��l� jY���
������� ��1��zΟi���8W_h��!C=�R��z�J\��� �J�'��������<Wf��:K/�|�z�æ�}�a��)��צ�?�1���(�1�@��3+��?�y70��9�"��QUf��`8�������o�dbS������E��;���ʳ&���*tg'�?21��X�rp\I�wkMW���6K�T96��f�y�����b���^_@�|�{�L׶�ѬDqtM���EcV��{~��`��g~��y�Һ3`����J�-��`hq�Hc��]UnMI����^�U��VpïP/Q*����4��mT��;�� �枸,>�#���� �w��G�6�)g�?����IP�
�<@V�7�$�@#S��Nwֲ��Zm(�1&�^&3�LT��F��:�i!��p_i��������j�Q�)���)��W��y�e�^����t�\ga~,#o�h�Y!��Y#�|ǃ=L�N��b�X��T���b��G��L���ɍ}t^ep,���T�t �'�V�w��s�S����(�n�a��OV��f��ϭ
���e�\a֩@��W��q��!;�	b1i%'Bx.\��*�`���� �h�XQt��K=djR$�­&x.���	p����߸u�:�n�L�ψD<W"qP��S��\�z%� /�?d�@Let�:��rP鮌/M�d;���u����{���#�Ш`�#C��~�ώ����Hs]Afʰ�����h�1c��5:C���Q+�*A��M�Ñ-:�B�\\*�&n��'w3%9�%%h`_}���tF&'+Q\��=ܓ����4s��O��PTE�J�w�R�H	mx������a�\���Ջ��[�t�;a48�C�X]W�һJӯ{�ѹ����G�c��2��3%[S�=ӫ�}�^=i�N�24�e�7�S���wE.�m�ė��u���~�̯�Ѓ�x`�bSխ�M���X88�����y�H�/@�15D���M�+�����?I��c���ѵ��`��#nY��ڜ�L7�fi�,ǧ���q�jF�z-&��_��')A0{�ݖ2v�A�#ӟ��=��Cx���7�7�F�6NBm��&��nec����X)������r�)ߟ�$e�Zc�; ��?������s1� 3�1�e�����9������h��m�3��u�*�n�c�mʬ��[�F�|��lÐ�fجV���L'�,;!�F���=/�G�r�̼b7���mF�H��
P�:��Ɇw��m�2e	�����e_�f'0�6S�����l�Ț�k²OBb�-�,X�)�X�^y�c5͂�V6�^�<:Ne��q�p�CH4OΣ�&`})}��S�*e�G�#�h�g����؀��ס]��e����E���I����k�Pu��>�,>�HĢ;���u�^��#"x�X���S���OF��a�|�"���d<�D߰r��\)1�+j��;���4��{��ȊE���m<ǩj�4����C`hd��H=8��Yt�9�fYƁ�6O{�y�O�|�Ⴏ�����4�@�GqE
�\<��7�MW�-Aۍ@�Q�W�qID��;˚�+l�Yホ\)r�_8��μ��j%�L��Z��
��'A��W��AY�Y����U����MN���륽��l@t�o�B�Yc��м�� ��.u��b�kC�=`)!׸n����Ԟ�S[u�e*�?�lT��765Z�hw�	V�wP訵���D�BaV��T!�D5�E,�*}#�

�Z��Ӏ���7��ů�wvZC/^� 5ѝ}�T���T���!a�U��X��\̱�R����T�7����V,���y8�"�[V�)���b|T9�lw��V�nA����|2�93�V�7e�ߛ4c�U�`�8Öx���u0]��g��ɴ]�`�w'x�g�����S�-C1�X�h��Hh1`*�����ˣ���ޝ�z�;�Fb�)(D���h�b��$�h'�{�I�6�%��1�s�<��aE`�"���s���]P�cP<|/ys��k���A;�(���GE2����}Ca+L9z�
C�E��~	k�h)�z�pk{1$�����T�Nع��g�mvܭ�<��X[r�V�'�zt����h�e?R��u��叿�Ϸ]*�O^�L35��G(�S�����RG�Ǟ5�s�=*�������t�"��x�0+�f=�s���a���R����HM^Q�F�-����6
���V�\���O����Pd�~J�WM�Ȫ�W!�|"�����Җ����k3ƶ�u[��ݫ,J`֝���H�1�A�S�U���/��'�s]��'�W�O�����.	r�0�cd��@Ԕ���@�诽+�q!�ou�ac�IӑZ�m���Cg�u�wS�0�جT#@���",Х8�%>�$C��=���G�q��@T2��������ʗ���d+�&�"(����rO`�>9�O۝U�
�á��x:_폴� ��Vq��o�l��g2��6�,��NlKNM��'�5��_Əm�A��)V�~$(s��cS��H{�z~� Vُ�^«�)]C�>9����~��t�M�IF��f1<D �fpL��8������JQ=�ɴ��p7�����}	�q�2�7C�!6'b�|RS(	��<��",��qT��U<�T�!����l�p4��,�7�l�&Q�͟��Ix�lȜ���ce{~V�w�Yx�4�LP�}�L��U�����Ĕ����&X8u�1�GU����3=��!�E��V��@l�a?^s�Z`��;T��"�K�:������؜%*j�^d�n�w���Q-��}<Ȓ/�F�I�����\��`F�IlԘ	�0i��==4�k`���\t^��N3X0y��{4l3�u�\�V�CtJ�6�Es�A�W%�G���8�Y=D�gI�^&��"���^v�F�ږ���pT�	�u5 �|82]D��d�K#�Mğ,�&�[*�mWױ�Q��f$n���y@g�����D��_Ql_a���4f�j�&�S�����Y���Y���4�ה93���,v����#jC�qf�9v����ڈUNנ2X,��Ke��\��C�������1�`>�}�L߱"E�P�w:߸��3g�up�	�̸�����ݛ«V1d���A��7D��$u�S�E���I�|t׵ �������{��~��(s	��1-Z��������IV���a�禱�� &fF �([�g4t��Az]��B�d��ږ�) Ǧ�<��ċ���"Gj�K����nB�W��c_��:b`*�b7�~�X_X]���ݕ��غ>@j�Y��k$���VEb��&p �L�%N��u��<�|�/��D�����0��?'W0\8�z������7o���#�<�T�şBl�x���Eq²ҷ���o��+n�,�RM-rݷ*�ъd*۵M�x撆ES> D�4Wb���:|�Ш�^��~d�K�sV\\������&&'CY1�][�J�����x�)?vd%��|��
t[j>Kۭ��9
��w5��?�%%0�f��O�1��=L��5�BG�Ǚ^� (׾2x"�Wkơ�֐���j�C�p,3_�^��]�8pe<#
����.�s}����U�{�!��C�K�� �Hir�b���e�ɯm}��g�C�?���y���`�Æ>�\x��)�r�\)S��������=dH^_�8�^�`to�T`�E�m���
Vh�m��[�v���D�h�Z�%C'�ׯ����zc�xk���m���h�$�4!�\nH�D�[,��BIy�P���[nw����`���1�o��n-aoRe&���VƢ�kܾ�V�!��Sv�IWZΨ�J���OЛ5}�bqo�RD�$���[�Z�ml���N������T8�Ѻց�V��yj@��l�w��1N��0'�;�(Y����k�4�����8sXLj�d��0#�QR(~�bUk/�%��0���o�O�z���͹㺢T��� KC۩`�
\wi�E��?á��c>/�n��Y�V,=4��Ki_�����f# 4~�}��/QhS�0E �<8�S�/��4ݴI�W%q؃�[�����O�Y��+�������.�����3_tp.�Vnͻ���5̫����XCg���o�|o�<]���h�F�B������S����Y��u:������L���3RJ�/���0�k���!. 8k�.�HP�
J='8�ü�û@ @���N�P+���4H���o�pQ�n/i\�\�:� ��^������4�U�`Q�X�nǲ�����P���jӉ����H.�!��2�_�A������|��6doJ&8�d
���6.0W����bi!��{s��
��E���G*�¨��W�ۀ!�CS>Ax�.�A��C�Q�H>H�i�m��H(�HQ� ���%��Ę�&I�5�bG�#͈F|ɢ�Q���l��I�����#�4y+�B�Y4o6~��'@ib���F�4V��~����2+ĉ���T;�w��J�m�3�͔ڵl���Ib#U�:���Rp���2?�N�� �7~��N�G�����t_L�7���������W��� �'�5`;���~�@������$)N�\���]u��s�:Pa.��cq��X��p���1Z|���'�=�<���Q���u~�P�L����K�\-�2��X�*�"�5�z��5C�����l�;K�ҷ�KaW�#D���wm�Ed	�*����O0M����E���m���z"�8.���Z5����t��}�k?���J��v���v6ȯо�����u{&�������1��:P�9,�[���B��ڗ��Nvt�s`&@�� �_6aʕ�a#�q��p�Fx�eݣ��f��<���D���ǡ�+�'�E�}�-3| ʊh0ܿ{��Ʋ\�d���M�+�eH���[��ָ�^�j�Ef��]��j��¦�{�&ӱ��C]ؔ�K���Ȗ���_���K\9�!\���f<K�o��2��y�ᦺM���ʇ���R����o�%��_��2�5�/`Z��'���+���Ũ�_�3v��D)2Ѣ��;�ة5�[�AԤ7��z���<S�jFM
� ɖ�q�b�]i���>������N��k�Z��X���6��L�Ǉ��͠}�w���]��ˌz�M-���c f,pzk�}�������~����yٗ蚸#��6Ps�Ѯ^�Q�C8 �v#��y/j�Kx����r����h7�r/+]>V���g;v�MJ�t�
T$�ք�-�����[Õ�˷ഹ� %�2
fo�6����i�+mw#Q�����g���H6	�b柍�Гr�#Q��K������1wI�״j��gK��fj�.a_vG�I��i(M�&� aCJ2Z�Ci�.���+�n<a�EJ�E��O��
[2N������ǭ�g�f�M�"� �a�e&�bN�� �ᓘe�����hrX,z��P9�Nx1��~nf[,��Kq7��lR�����X4�G�H:/d~>)�4oF��;�Q;r�S~SE�kӤ��'���"���]������)W�H�LA�mc�R���Cc'{&�w�d��ޠl���Sro�K3�]�(�0��(0���W콕�";
���di��o����F��>Z��,x�r�����;Rb��Er��px�u7v��l�~�Fn�;AD��×?���ε�?�kX����|埍�(����ju,Jv�u{�To��%2�����N��kx�l�b���ehl48�GNx�����$�)�?í��YL�Ts�ɹ��Ǒl%ous̺Śځ�g�K]�).���/�w5Y��������Ӿ����J����vet�	�Q-w�v�����C^b��^|-2�|T���ݝ�ܪ���,u17�b���o>��^5��/�g�� ������ª�x���je�!�xEk�m��I�:��
�e��p�����;'J��	6�F���m9��D�h�!E���b答�ׂ�<�Vד���<���R�'�2|����1m���T����1���9�f(�G=88BJ|\�If��{Ӗ��Q7(brR����1ibQ�����Ճ���� 5�f������*8��/���Uv'.�}�w;RC�Hm��N�>&ǽm�A~hfF�is7h!��� R�
�+V%�6 ��\6d%�;�6�7y����c����wX�@�*���9��	d���6 ��3e¹.�ڎ`���!F�<9�E��Yv��?1-/><@y�^,�����p�b�TW�^�w�K2�ZP�%i�ի,��+�[_���."?D\C�MTӒ�]��S�۩��@J*�����g��øHBOD8Hw�^Zuј�Nj�RPr:a�4V�����{i�_Z��n�'��D"`Dr�߇I�b!d(н8�Q���3�C^8���	�?�(�!�K�MǧH�r9ʟ�!/�1�EJ��MPq��Gb��♦��˧_u����dˤ.--�@׀�ܡ6�繧�-F����P�L��鞾}r�V�ʍ�oG�D)�+*A}98���S���-tq웒�n�܃��h[^~�^E]5�[�eTDR�[��0����NI��a|��荩�����gWU��Rʄ�{U����V�����^��RiS�70`��p�e�C��f��12N�wc���5H�O��u�7ھ��8q��C�Rc�ȭ�n��� �?4���(,��`�?�ZJ	y���'ͽ⧟�q��]?��|J�b�.ד�j��)!�Np�)R����ib~qOJ�N��te� &��<����C"R�C.����e�:����_
�9@���
 �U���1W���oT;ƧH0�Q�����(w	�ii4v�M� �=�R{}�\�?:aɠ��5��L���}WC�aaE���|�z�ņ���`)�ʹ�G�Gg&�h��6-Q�� m��B������k�m�>/b4�Ͳ��ZU:S^H?]}@�U%xfZ�|tYJ@tl�J�*|�g��Z���o�R%eiF���B��?O�6 e��jJ�Ψs��F�i�=\,�����j� �5�9DÃ�9��wjcL����Q�X�@8�cSt~X����ɘ���l]���#� ��q
/�{, ~��[1����A�x�1f���s����t �R
��p��<�cQ��CgrӡN��Npf"�8����(��!礒�q�� ]�ͩ��u�\D�<�Y�_7��A�X���q���}>��8
��[@��ラi0��@(L^��2��D-�96Fhw��� �Q�oI��ІN�I1������q�ѶhVO����'�y������
�#�zr-l�$��x�_�no˓�aD0X�,w�^�c]-u�y1��� V��i~�7���Wy�̅L�L����-1��R�E���7����g�KjߑSH�������<��i]�N��x}��~q#�m��럄ycIK��v���k,e�H�u&x��y����z�B��Z�%�<h���nHsI>�E��y6$�&96&�[k�м
�(mX~#����� �	9ǩ�$�bǺc��MR?7�~V]����Kي����9�]>�����S���B��S��n[�#����1,@�n��o�D[�G�$nGx��?�CC��**�Qr(�^�1q�����I��i
��x�-� C�#}ou[��2��Y\��{K��*Gc���<��|�4����)m�*���(9+���QW[����K��.I�ֆX[�'6������n<	$��������C�X�; � $%^\�n�C0��I��sb�ù�- di�w�8��HLX�!�?�I�����HM�p�n/����ǟ‧��am�>�9�����tAǟ}���:t��a���a�#��X�jo�b��l<�F-{V����Jl�Y��wn��]`Oh��Yt�u�}��x\�Qؿm�+}b���|��h=����y?P�M�sy��n��P�2�P���8��w�C0���8B5\U5~le�ޚ��#�_��&'����ɺ���W�����-�?����ߜ��"`JE��{����DH�4	��=������@A?�k���6vp��8po=���X��rO� ~It����(F�D�5@�rl�)�M����)G�5���B;�(e}�>�CǇ%d�a���"��CJKh��$��}�bZf��}M�� Q=����	 =�t�,jc֪�X�i�t�(Wqw��dMN=��^���"y�c��@j����k�x-|�F�5��s�ɆZ`Xzz���D����|�F�ش^�l���٥F�ڀ�HѨ�Sm2Г:������k�\���;���+���w�y���/�|��]�p��5u�V+ �9�Ye�.GT�q�zqK�h��d�t%���.�O�M&r���,b�m�<�e$�X�y�:��M;��蓵���ߤF$��1j ���'����9����!�9�}����e�,nէ�~}���G��J
8,�Gڈ�}�� A9��'bA0�hTam^���(�����k%�K�������u˕���4�BwPN^Y�ۡRV�A'똳/g���׹ٺS�%�tA��������TL�s��ڰ��ޕH�%Wo` ���-�>IJ
)�DI �m^h`X��W���,��̨s�ސ�(��( 9���Q�Ju[2�6I#��H�9E���u�B��d�=��3߄@\���+c���>�����mf�)������QECYor��j��΀��j0Æ>�@�4�*.�:,�v�x:V8Mck��+��R-�sO�8:߾,�Q�_ZH�� �.��U�|HM�;�L���]�j�R��<�N�_Hp���e*�+-^iz2�S[\���-�$X&����;Ҧ��Z����bp�Q�}vg �O��4�;�<Vb�;��d}��:�lc���M����A�k�zRP!��������	s�{&=��s�[�9�eC�g2�FRO�y�խɕ,<r�#�G�c�MT>q�'��ok�w��p+��>ޏ�+b�܋E[�BpH�)�>���;!T��M찍[��������ֆ��>��w|��0'1sa3A�C��hcTqL�+��}���Ek?8d��sCh�5�N��ޚN�V��37|-j������Z����>:=6k/:��˰���@@��}\��c�1��wٖy~g�� #ڽ�MT�	Hr�=��wb�ˢ� �@	�+2*���U�%4�b+<�(~�" ��/�Bf�D�`�n�|���{\?����	��P�[M�xr��d���Z�c�5��R�Չ�f��t@�!��ɘ�/����#ԛD���Is!�9w��Z�f���:bX�}U̕�V��2,-�j�F������!�O�eҕx��ѶPxem�"C
�,�((bX�be7FW���'W�Hj�+����7/����n*|��͘=ܰ��Pn=lt$|�M�浓CrO���&�硇�B�ﺡ��Xk�9�&aݸ� ^�^�����*����I��=���R8A��7�W}짓�:���I:[��A_Z��=��c%�8kA�4̠KrB���	=�_��;��j��[�K�d:˷)%mE��W�r�3������7�S�+Ծ	����5�/I�7�M�����S���4��O�SH�������};�1\-�1Ɋ���"`�a��"����A�S�s��$<>sJЮ����u��]�f���[��fn@EƑ˶��\?�뾙�0��mL���&��p`�yDͅ�R&��c�oQ��?S��_����Dϕ�z/�kl�
�I��/�􄧭q)ȨH�}S�Q4.d�+�J=��V���lO�\A�<�w�υD���_Vp���Ż��ܽZ�Q�.¡�b�rU��u�Z����O�|�m4��k� ʋ=X��o�xUN+U
��?`���J�����ut����*�:F�j6�>�������)���#����֖I�Wc7�!�u1����E����H:G�8OW]�ͳ�v�	�Zc��XF���Tϭ��a��Iۡ���?�UZ���tof!x�7�rF�Ť�OU\��B_��ߔ�ܷ�����@���^�g����>�69s����\����6A��36����˻({��$D����?"VbYCJQ�%�f3��7a
�f���Az�֚���g�^w4@�;�,��9���YP���!a"y{*U����r��ob�)	BMc���O�)�P�:�/&F�7o��g�4G���)��+�P�X��~]P>��ul�\#�u-<�-�)ih>#a�6��:D����0I��$E~JR|����c�5�4�����䢕ᜱ���G��íz��7?��l��` �3�X��K���_����6	���W�h����w��~�f�q�,�J�n����)@�lW��P�!���lz�F�[�&�E��`1���Y/u�0RB不N'n͙�呝"��$5�d�s̸�t�y�u��v  |���7����r�>�-�T��]�Ϩu3!�l\�t�wQց	34�imP� /�Q�ld�W#7û��C.�zhr8�ǿ�}�������E��1��8!K���JE`�MV_�u.�G�I ��@��2�@��j��s��,F7e�}$�8��m<O�e�ONO���,���Rz��f?�Z�\�<&ߩ:vD(�M�+��[�S��N�r��g�n��C����z!�7J]Cz�:�����)l^s���@ؓq*Xhc��t�-�ւl��▤�d�>�,���$�y>�oef	^8��0V���[��O�.��bg�8��Dn��D��/�F(fj�=�x�H�����S�\hN�H�:Q{4A�,�syrSl�p��
W�����x��~��pY�+b�|�o�4 �PE����GlK���+���&�9���,�
�`V��YπQ�
��?�P�û�x��,>TH�cu��(p��o>��@������3��p�_�v�Q�b��NDO*xWe�'��Rc�T��^���dnwS׬?�$V6O��o~�u�Jܘ�]�ϴ��z�p\����uX�L�����Wb�㡞nQhK�|��.,cŷ����g��$d�-�$�D���D���5Y ���R6L�	���?�?1�p¿�{��9�S�%(j�E��$���x�w�_�>(#��7a`lvYԛ�/3�6��"��1s���H����8'�9G�M� ���x����[�O��+1?�;�a�|	~��)�[ @�-ˀy͋&͒�G.>p#H�f�Ĩ�#�P��꬀������=d�l���g���\'�f>�+{�K=�5'�	"K�b�ǫP���\��CpH�S?���0*`��U�<�����k穀D�j���Lsn��&��{^��c�,7o���gA_�Fsj�ɞ^cs�^���@�dd�k���v\�F�Z[U�w�j6���(w.Hf>l��SxT3���n�������
�]J$ve8��.X�̰)G�$��3i�_K2eG�E��R�#�:���/`�S�S������a��m>��x��0��L��u�m�Wo��4���Ugij����W�Mf�U�AX����Z���Q�|0Ɛ�ȅޗd���&� =�H�j����0U�)�/��gJ������rZ u�Β�	�xF0x�7?��,%�`�K�e'��bB�ϰ�XIЃ�O�Z)K$��5�^E74^ڞ���f۽>߬'J�\������g�>����o>_l����s�h�(�Zo��^Ј�ؗO�ڊ�����8����vљ�n:6��jݚpGu�S� e���oE�������)�M�a��*clɀ�o"��������c�.P�=�%��1���3U�<����^���F�N�>)���V�:�E����?+\���{�ǧ[�e�G���W�K��:Y�q}yȀP ����W�%F��u�.:��CR���I��O��{JY���g�fP����F����r������Lkv�&(�"X�5w��:rT$}֝b���UL,�H��`|�� e}rU�2@�����	�^/B��<8�	N{�������!�5��d9y⵮H�U��-a�7*V�7�%W������y�M�vrC�F�ߕtq��D��98ύ
*OAd�\D*G���o��B�L'.t�ط���[�Q<. Y2�~��S��4��<0��u/=؞�2|6��{E��G�`����E�"�BZ���C��:��#�inM�uc��� ��8�ws��ݻ��i3!q�6��c&1���i&|6D HRJ������W��b�R����@0���S@U���C��^�F^#�LBQ��=�{iO�@�ҡ�D��b�2g�� ��׺�2Gi�M�0��ց)׿CE��cc\�I��D�d��0p�U���Jc�oehȍ��o譂��yC|���#a��h/EuX�n|��y׺��bq�m'Q��X�U��9�V�
}#�P�3ZO�~i3�g*4�驋���ZtX���i̛tuz�E$�XS��L����"�\�h\_2� PͰǵ5�H�N!��aLH�$$~�E���7_�O��$�îg��/�O��;�s9�0�|�Sⴆ6.�������o���#�dMA'J���gGy�g����n;?0�-��`u�i|�-g�"�4�5�/=Xp�)z9�~��=�E��|Y�Hj�$�d��|�2@��+�R~����^�aW�9��>TN���
iX�� ����	��%i>�3O�bB��hV�F!r�t�^�b~R4�8m��ǏҾ����J*�eN
�0���@1'�7�U�Qk���C���N���,�9�B��_/Ma�2�q1��7�����d��uCЊGc�X�_U'�N)j�>7L��
B�R,sI^L�ea�YB�&;�Iv�d­�t̳8� �3S��*duO�����v���3�����������\��~� X��]�Ŏx�S0PO�G	�� �KwΧ�=~Yy^9��4�01��;�D�S9���]v ��pB��&ͳ^�^]����C����#��6�D���!�.TA�)�:����ڰ�I�kF���G�R���Ǖɠ�*L(��Im�&��:�]��(	W�(��˄1Ρcx	 ����ٰnH�����g����v6�!�p�G=��Ki`��͛��v�*����F	!������j��i�m]�+ /��z�2�U[�x��Mv$��\_'m�%Cߺ��a�����/1��-�f���|��։���듆�ŉ/3O"�ݝjُ�y� �V����� ��Y̾בP�Ġ�?cGA��UZ�q*��o����,���t������>��
#y�)�q!1v�W1��w�G|#��S%�'t�4E�Q�5EA�k�%Q��+,Z!ނe
?1aY��#iTW��+��y#σ�Ts��E�Q���q,\�_���D�����r�mBv�}��
�w�n�X�{�S?j^XxH��Qָ��V�(��{Y�:keƀ+\b���\��O����9���j!ɶ��!��e��|��'D�F�Ub�+d�2&����uK�9e~��J�2���;RZ=K���VňJZUyi��߿�J����Z�S�����_-y�;Ef
� E�"i���{�"sF}]�K�T�1�X�,�T?���(S:�tE��b�2]k�c�d��0�@�P��h�]]J��;�~��T��h(D����8j+��f����m�֦r���q�Cx�[7��/���'�,'��t|>W�aT��na�i���{bޫ�c��BrL0_����L����1���Ӽ2M?�aR�v��"_,�D��5���B�J��t9���"��U��� ���7��e��E3©��<<�e�U�,j,l'�eQk�h}jY/�HU��̢��\���S�KP!}�\h����н~��C���8�6�b���~��C�ʸ���fo>�/
���@
5|Q�ˮd�y�`��!������{�Ng��r,~�����YX=��&�L5�ZN�L��H�D��e<;E�* ���?�x\���xP�:�j�[ʹ7�<�!;!��YG"Ɋ���J��S�*�Q��[�r�]��ӮTu!��������+T7b@�T)��Xn4�倈�ʐd߃�c<���Og����B�%���u�Z]j�L	���?kƤ���0���b�Y(�l�m����[���D�fr�*�sUn|��9��n���{�W@���0��s�y��o��b�UG��cxtp�~(�rL�ɱ��mo�4�^C�&是�ײ�����)�+�yn���+��&t�W�Ѽ
�VD��7�M��`��,8�!����`�~]��\�dT+Rf�S�_�+�xۼj?�
�O����|4�o�lq���{�ͫ���_b��1�Ɯ����X�����W~Y66 \/}>�7-!Y%�U� uW�T��	�	C��ڔ�a�ɏWc��l���â�Y�J������ �_���D���y�"�AvD�dͧ�\��m�*�RQ*F�ܘ���J&>���G�e7�:��.�Ynhƺ\(��)q˵��J�	��H:
f\�� �E���S�f����g⛏j+)e���;�������|�]�JH�e�h����e�|5���9�h��!��x%N��O��=V�<��*���cp57la���|I1<��]^&$�iٺc�ڹ��-z(i�t�Y�l��(��o��͞�����D�^���"����?4G��_('A��_6k�& a�w�^����rJ�Ҩ9X�쌇-\�q�w���v/YpK$ֺ�C�d�����fQ�I��ҋu�m�t��������!��CgJ=A���rȊȺ�`J�^ZOv�C;O,��^�]��w�!nw{ݑ}[�c�2`0�"
{Q��_	޶���ڐ�T���������S]5��ji��q.T%a��ٜ
��Y�̡����5�0������h�x��\�g��>�xB��`Ii���SXF�U;��Ε��:�`��O�t��A�M�k��Xb-�sӟ��Z9T�3`h��P+�|8��P��E�3j(��I�E��Gw7�����a���Y�-#�7 \��px�+�Q�^]�S�^^\?���_R���@���!_��;�޽j�ە���� 0�Ү7��`I0'5�Z���Ms�B�F���|�ς&)��Ц)��_�ש�+ J�:��I�N"qq�4���T1�д�g��g�a��Do��D��r~-.(v��[H�� ڲ�� ����9�������.��ܝX�t%c';�F��A���u
,wCyg>��"^'���YU<گ�A
CE۳�Z`�⪢J�e%� jOV���Y�7��Mf�`$ٵc�a�q��q˫J0_{��J{7�̧��λ�ɩ�~��ĵ�T�;�����V\�Ig��	b�f�<>���/M8vt37)0�x2v����;�,�Sၻp�U�v��$�7��b
w����9/�
i�Y9G���D��j��p�J�j	+0�Jdwl����|�2���h�d/8����+���o��d���&s��F�����1[�X� B*���{�q5�{��Q���*���W{���	jcCHv������[�=S�YQWQ�����mQ��6 r�U���;+��_�|Et�V�ZS�H�%�<̥�4�a����B�-��芕�2k=�]
B,�j�7�ڂ�AEI��m�u8��z�,��Z*4Ϊx7�E�`�&�E2�ĝz�8�Àr�-W��8̹�M���̘s�g�;��$�mϓ$h��N!1��ԍ�?�0�N��7�Q~Ϩ�o��o���8��5L^	����BZđ�b���ֵEx���k"Y~J���XS[|?�i}O�U�r��8������4�8���K��l��V���[��Ww��]��+�f�����#��ﭐ�h% ��kᡍ�Ԧ��a��ߙj0��h�*�A�-�肒�jd����
p�k;Mi�H|0O�b�����y� ���7O�]G�1�-gl5��f�pv	��%�D���EqW(�'{v�_��I#����v�B}�#��T1�
$�ۧ�y-�d.���q��#�Ǫ�|��GCd�eb��oހâD��(�C[๻�;��0����)�
�[#w���s��`���ߐj��n�!�d<��Ξ��Ey13ע���B��Ɇl}��el���W������/���[b[}����ZH��I�1s�%B�������y�Ӎ�L#x���#�)G�����K�)�q���V��,J�������GW2l/��}�To��֐�g�Z<�R�EL�(�|�j"a�����K+�*�R/	��]{��xt��@��`c���d��Ǹ��.3+�.ЏIM�F�M�TTi=+��B�yy�RE_�a��T�i9e`��m�Sˌ�79r�!e���-ȭK�:9�����Y�����y-����Q�lI�$)���/��H�p�,���)��X�Yd]`�N����1P��I�N�b	( �s������M�1��'���ة%�J����m�+gbĘ&��v�#���u�;�2����R�5ot������ T��l9V;�*�}���w	��-�џ;���0ɍ��x�nfTӌ&��b|jO������k����Vg�uM�����K����������G9us�h�����'ec��oVV���֊��Ҫ��MF3��{��[#�TN1�P�n~R�;�Лo������
O� >A+&ؔJ�\f��y�۾y�C��� hO*y]�υI"|��Â-��CN̓Y�l�L~��O��fw]����Z��@��d�(ˈ/��Ta_��Y`UD�x�v��E�Ӌ�}f�.�2 sM(9ðP���o2a�h[
�� s�|},�bQ\�A�p�vN�X�)�|�0���4 �jF���!L��R�$��R���Sѻ(bD��R�J�'-��Yѡ���j�ƣ�Y�@�NMY~e��΢g)�23D�9�U��ڂ��dj��'t�S��<���So���2uy<��f�V/#�=(���p1�nLϲ�uX��U�L�����Ɏ�{���eM�^~b�tqf�1�W�f*�C��� ���&d.$2��B�:X�nQQ�\�o�t����;���N6�_]�9��b�Xv���<�5#�_�Jp�5���N��٤�z�wP~j
\�Ƀ����J�J�y�S����#�'�����YP4�V6�9�N���:d�� }̨e������LL�飭k��9y)������VQ�W��/-2�m���H������������#��64�������g��U-����@%F��;�6����*�lݝG5��b��}1:<�҂��d�Η:D���U��e�l�v��Zx/pǨMa��ޡ7K8������Z��0�^��-�5T��W�6)�������5گ�1�Ө�|-���|�����0��Z�Z����P���#��	���2���r�,'L�>Ɂr���x��O%}米\�6E!��+7"h���I:,eX�2l�ך��>���/E��YnY|؞�x���.bzB��gl=;�$��B����gYU�o	S��J����i^�rk�僊��d꘻���-�7o�:�~
���8��_K���@9T�iSH��4����3��<1 �h����]����Ж6�cO�g�
�����G'IM�X��qq5�s����W@ɮ��S�؞<�Hk��^��L��$��+��_�!
u�����#�x���Bpu��,��8���3[�h;~B�\���z]�ݏ�O]�(�jͳ9�5wd�������Bϗ��v,��8��rT$���WlvF5%:���4x���KIN6?}��97@���צ�������9���9�.�=���w���k��j�E�������R�[,	�HB��n��yъ+.}����u�t���:��Ð��65%�|�K��r�7�u?���r�x�[nN-B"�J"�j�ip�s!���S���N���9Xk;ު^�3�G��v*�F�A�.��[ܦp����r����R�Q!�j�#��J�T�YEI=Ȗ���i��]��E��w�c�F�� a��A�ҋ�~`}��5p��%^�����$��'3"�
�q���-G[����s�6��i!M�������f���J�̎X`x���qtQ�O�r�!F�t��~���On���>#J{F����\�P��[�&P� -�B#�5��ǭ��=1i0:�CC�pv@[ŝ$�.�=��h��`�xG2?
��d�R��d��Aɤn���t�=Dx��p;���[���i]*�׿bu�m�8BS�z�� ��;��Zha!A�-Ϡ���9�Nu߀4�t�0,�>�MV����0h�9�]����'xw#vm��n��Pf��bƺ ���� z?�&�.L�L\�U�;�-/ޕ����ӈ�؇�O�
\�Xhk�[�g&{0Y{��ﲮ���e�����G�V�9^�7�"#�q��g)�A�Ž��=3N񶊥��4�4�)s S�*�����D'cЊ
�<.�ud?��"�����}��	%]���[����rȵ�`�����p&n��`H�ˤ����S]��.����+�I�Q�C�l}7R�F�
@ʐ���NU?�~ɥ�	$�7~���	p3�U�Z�nS��B�5^#�a��fq��9l��o3�B;����r�XJ���i�+��w?�V���I�Y W')�R)�8_,`{"OzI@!�-"�]����I�^/�����f�� $��Ө's�H����<��X|� �#:�<,V�������'� �5�A�)���	L�,�V�Nvظ&������U0V�N����W�]\��<��ujx�S�L��։�-m< F��XGM۝�y�ri��� �˸D����;	BD�*�,-X<�����
�>xY�d��U�/�7�� !��R�4��s���,���K.��d���o���q �w�]����<��v��s��]⫗�{QP���HR�[��@����d����C�h�&�����9!�ks��dߟQ>%燛U8[n�-���/
?�g~�����i<t�@kS[+�!�Hu�fq�ôn,�L/c���+o��'K�!�~��巖�n<�Vs�z�y��5����X���!+��s-�&��Ő�X�U ���-a�GN�m���Z�@�ڔ_���t!������q�Ә���֔=zSf���8G"p�T�<	�.���;F΃֞I�8�Ң���`X��l�eD[r8�O�c��>��Z�ߞ��y���&5�#�L�-%�u�˷�mnem�]9��Hl�.�7�L���C���f��*�>�IkI�E�SP[�Ѭ�a�X�qRr\�$�o� �1��˩�<U< ?�������X�`��JC����%��Q�f7Y�G��-YrCbht�PmO0yC!r�'\�a�Lt5�8Ve<��)՟��J��<��S�/�e���>@eN���k�Hp�~�;^���Q����2������E]��4/�ԯ�QB����g	=���-�C�����RGoQ��C�]&pS�9���F���=,,�0d�]��7������(�DK���l>w6�w֠�I Sׂ�P|]`��w��=
F�pa�ہ8���LY����q����zļ�T��VV���m�i�^��Uq������M@�<_RBBk~�灞d��ʠ�Pr}O�M�q���
87oPE�8V�hm��>����ML=1�`rZ�.x)^�H��^�0mp�P���V0�~�:%�6�D����p1sWF�]�9��Ӧ����ˇ[U�D�=���dIS�$���\�©���
>/�7BRr���P��U�����
!�]
�9�ڲC$�@�x?�]��t�Ol�F�����ڱC���G���
��q���bT��D�jz���W���Ġn��h"�v��b��ao��d�"Ȟ��n�zy�B�4A�-��4d�.x>����2��RƗX"�AՍx���kR�s��P������[j���� ������
�����l	������������~���X�\�9�+�S���,��h»E00��``?LR�CX��ʂ�>�$�.��y6w���wrk�zJ\��n|O�@��YX�����v�	NJ� g" n�B`��t:7~�����A�3}�i��}k~�?.<mH�s�%��-CM
wڶb��W"�쨌�n}�#�
 z�+����|#Cîtv�ˎ�n�����'�|��o}�2~E�p�J�j�g�\�ۀm���'�@a�z����Q�v��X�f�L��(U^nƇ_�p2bL�4ޤ����(9-���q���@�G�����(�,#���ۓk�"煮�����3�:�w�ƋX�w*B�Ǐ�X[,�(;uΡ����Kq�0�R���܉�Qt�c��3�^�4�7��ju�j���t'����tC^�Mt� SD� _�Ap1����0W�Ք(^�A��%Ͷ����$�
G��p�U�)'c��W���������k`�����*���'��k�s��k�)v��ЍV�$hVp�m�+M�UkXQ����O[��JM��7�b�F���K�u|?��:TP���C�F6h]�Q�(X���/�R���g�%T���1኿@3�Ii����ہ�#������G=3v̠4�~�W�
!��*kf��y����;1z|�u���vPt��v�gm�Mm�d����Lx������$����4S�{ˆݲ�5)M���Т_�/_C�b<� �"}������wz�e������׷�ɳ�SR /�����d� v�`��Kf}�NP�ު�.�9�q���^Ƌ{�d��֏R���Z����k�C�!c��#��z��6&g�mۦ�)mV�Q�~��&X}?+5V�no[f�Pv��$\\PaH�| H���n)|̬���Zy ��I�
a!P���Wc����ЎK���
��&�S�' EXk�����/P@�����M�}�pJ�x������q1G���ׁ��e��Q!}(m�`=a��l�|\�tb��;��Qyv�l_G㟱��)+����o<�����c�vv6e�/+������SL���:6L�Ri��(br�L���r��m-PoS�Ռ
����tKQ��\V?#Y�+8 �"�)֟27�?u�X,םK����c��0���G+Z���TH�U��a���u��/�!٭��t)6��_s'%��U��J�B/IOIe��dN�^�zlAA���!�T.b����8����gr�������=^��hS�@Ja�^w�by�Ԁ�@UP�B������i#����V��+��R�t�,2��ōL��yv8M?�"�+h{�6q�����f0���6M {���E�<��{���y��(�d�l�$��\�K�"o�	��<��a�OC��I6�<�-d�b�S+��家{�Ǭ�SCT���� �IP�մ�$~:)A���?4X��4+��;u��>:�{M6�]�M���#������}��,9�b/!+�B�w���&c�P�4��O��]��)JG@b����/w�m�_��A��X�*�LDѴ�yH�C����,�����7�boZ���FW�������.>�#Ine�3�X��v:`�a�˳�ˡoZQt$�!�ͦr�\������S2���C#SD���� ��'�T�4��8���,F��w/�;�_�����{>h�g��_�N�L�}X9U�5y�� �q]CW%���r�G��9d]L������cǭɘ��,c�Td[��墀�E���ȑ��h�W��n�`��}FZ��M<ژ���9s8�� ⾚���]kV��V֕�f��s)�uO�KQ��>���nԤ�)��5��������w���(F���75`��,KQ���@�lh�,J�¤���g���7��6D�l�g[G���
̼��ebY�iL��]f��4���st1rF���Ӻ^*�$��-��"��.�Q&x�7|�J�l�B���`3�<����}�h�;mS6�XR]�-��MNuҰ7m����U_<�ҕC�6�2;2�=<�ʑ��qP�᳗���Vs������N9�|q��Y��쵕��8#*�F7�oB����|8p$2(�ؘ����r�+�X,B��l ,�wL9Y��eMS�ɜ���!0�7����>�a����$�ŏHm��VS\~�@��;hg�my=/�;�F�i�|jt�;4aNT�T�����'Z\�~8��:X�P��6H�Yc�b�|bS;T�n�I�NY�wa:��X�&�q
ᑑA�����(�'M�ӛ��ֿP�@���q��0�s�B�h�P��+����(�����ݝB�)�#�m�M,�@Fоӿ�?s���e&5�f(�H2�r�z__��wV+���O9�}��Q^i�dƲ��>na���L����K0��;���]�����k�F_�K�K��,)
.�ҕBJu��\��ͻ�F��edq+�*G�'�v�d�4O[j���eD�'���mH���P��H!1��C�r�O��At��� �VExY6�o!��<y�%j�c�$���j4�$5���cE�Y8�s�lx����LhS<����Y�������h��������,NxT��skGhD���Ω�O��(�����`�t�5_t�u!I�o����J4:�W�ǋ�p)������O�P�l:/e��~��#N��䦼@�M��{���Lё#ݎ�~��B0U6�]��zR^��g�y��N�ܠ���ݴ|�G�^W���ygO?�jCA�GO��ɣ:��w�	���#���;�Nl|n�	T����I�;��¿'�*�Fh)k�y/���N`��}�uz��G�@��i�%�}�<��Ʃ��PUUC��Y*��Yf1Ԟ�I����Εi�N'�#�"c�����s ����-o ��F��7HM4���0A�ڿ��N���4K}`�y��UN�hC1��G�����R0�� I�*69��KO>���U����Ǔ�b�қ�?F�#���!
Og�EH�SA�6�eЁ�*1X(���\e���C�^ӻI^���n�{�cx�S;vpyˡ��.�^Y´^�f�)��8>iG�4Я��݄��P�f2|N�_v�C��_�����hIr�i�͘t����2gZ��Y���"�E�Ȋ�\�؁��� ��SG�� K���v�C���y&��Vx�Te�B��&�h�B���Vcr��ĄQH�׼�*����B����'K51r�VE3 fK���-�9U;���0��EHm�N��Q���X�˻ 5�#��ʋMU�N[N���|L(p��6���f��l��g~G�z�,Ԧ�X1(�G&�Di���ttz+>��|��-u�aW�j��4�Z����l��V�� �M&��F�L��N%�I$���o��Mso�~7��Ir�
i��0����=0��.'C8�š6�Ԧ'9� �2f,I�l����4��z�إ���ظ����l9�%qXx�����ë��Q��io���k�Ӗ�ǂ��L�y�7K�����+W�5=Q�Cc���d�6��y͜^}�%���.�;�;7�a�H�/�������Q��9I�{��\��o�[)�a3G�5V��gm<��/�C!O�ƃ��_��S�ʘ8��M�<��{��Fﲟ�.��C��A�]�%w��
�0�.���M�"�k�;��0eN���b��Z���*%�
zbͯL��t)���L�����3�ŴM������6flj��XCG�j��-�f��SI~�Ğs��۱�fU�]300Y���nS;:�_��@�$��M�������!��%c� [������/	���DM��gq���ђ��P7�I�P���v�L�O��.b�(��w v{�`w���/���X�jm��y����)�����A~�0��B�T���z~a�� \A8 No~7?{��8��L�k�z�~�;����/w���(����q�!e]���=�_����Qa�K�L�C3������i�N��L��ʵ/c@zH��Kg5Qш+�I�V|�"V�J�ǀaO4u�$�`��E��|䱿��P�����#kkjZ%Lv^���N��^n�LC�9s�E�ο���W~�y�'��4��bwpS[O�����-���H!�m͏�X��/���#!
Q!Fԓ�1^k䊝�+?\����Zң%Ǵ�'X��'ǯ�3#"�����q�t1��8�V&QD ���d3�La�(���:�Q�ɡ���b��0jn,�=P����2���-D�9���G�Z�A�v���Y��7	:Fqv�Ef�5F#�߁A����\���g��}�R�DY=D7S�����iBOi�I���顨
�w[�6���*	����I6�oħ�
=Q�2����P�ȡG<�[&���,�&'�]�ʰ�_��� !/���s��e��8�,���f��������%g�ä��o�P�RF����5]��U�׺�e����r�v-����}\!�a1�_�(�OEP�9��Nc�M'a�Β��mm��e e�vSuC<mY������Xe
�4N�~J:�_�"ɫk�����ML�0�%
@R��Q0}�ʻ���l*�$5"D${��3+3?P��se�NRщH1"y��0��{�R��V�=���	>|&�?ۦ���ȩ�Ʋ��,}?�����矣�f�I(qh���v�d7=��=mՄ�ʡ�����3�}Ѽ"sѷ�r��� y![�T"dd��+��mX�E�0	*G.�>�V
���E��?�%�fH�_ <�ʷ��s�nw�7�Jه�v�;]����{�f��;U��2gRt����)���."8��m������vr}�j��Gҹ�B�Õi/k�)���dJ۵�9�
y7���	]�$���JG#�}����/�0^�
B�x�;�?��Ҹ|V' Fh�=G5߫��"�Zu��UvW����D
F3�O��M�x� ��%���0���P�f�'3v�	:�����9
,]�P���8%���>���:����ꡦ��s�uX�1٪�Tj!o��u+w��������e�oZ*���~*NC�@��H��F{���7��mT�
�,LG���Dm�g�����������W⹌��1��n�Qq����-��f�No�VY+E,<&��L�e��*U�E����`��3@��P�y�w�г>Lb��|���MD�^�ޞ�?���]J��e���)0�<���#T_�'��i�8��UG'�B��w	|��_�ːuD?h?I/rK�o�ό ��Hm!�#T��&��_'��k�89A�ERI��T�1����nq������/���7Jo0�Y����>b��6(�7�8Ik1G~�V#���c��*P*X%0�"��,)J��1b
*����5�(�~�_'�O�$W:dy" kysC["~��uq��#��J�Hɨ����l�lB���-�j$$>��A?�=�.�t�;I��s6ů��C�]����	j��kQ(~������K��cC�*GS�i��$�S)Et���e0�G0@�E�(�q��q���D��x""��dčف_�.��jc��YmCt�~�$꘠t�2�^?���٧�:g ,zy2����h]�F�C�P ���Q�i��w�Y�=����ޘQ���ժ����8�?��)[��p7"� ����Wf:�d@C���
LG�S!�P���8���ή��E�|�����t������_�C�x��zD�L�J�~��!E��9h�SyQh:��'T�,�!�'J���iQ ����L<\�׼h�*rw��V��$�a��y�.2-;�ݗ;d�������4=�_��֛5�RO�&D��5��F�bΚ���Qx[�@Η�)k���x�{��,�Q&���l�["�"�Ê	�����&S��Sq��r�`~��Ƹi�
��v�[�\��W�T�	
�R��Z�X�`;�	�1��6*I�5����P����-Z-���!6B�R+|��@|6*��u'�'8��	��3����0m�Ѩ���V�ɉa�:61��t2P9�!�m��&��8����ٷ;�Si�:v�9��4�!}�(8*ˌ���y*�f�)�q��3�*����`tu�����|��W������$���ݸ{w�O�pJX!�ZY&�o�C�u�c�����`�?H��U�\d���:\�]!���'�?�q�G�>�f�z��wԨ�y��F�l�#;�{���E�?Ir7�	M����,B�7"y�sʜ;%�8�1d���l��R�Y�z7k�4�/���.+�[N��� d���FM�KB�.��)�/�|OƄD]�(��krQ�flBD�,^�,߁�M#�JOuC0�;������r���>�>�uSH��k�r8D5�u�w'v�;l/K+I��>�)c�œ"��L�g�o���åՊ��2�?"��RF��ns����m�/XAz��Q-t��5��׆(Q���ܠ�Z�\��ޅ=%~���D�}*���͇g��qke?!�����f���������Z$>	4�SZ���S�@���x������M"9�c��g������%���}>{b��8�c���k�JƬ`����'<a�DE'�4���͐�f�-)%i��~��pC�J鍥�H���0T��l�U��]�l��w���#sGe���M�O�Å(e�i���o3`q�B##xM֊��W9�R$�\!$���X�X���wO�|g~�+��{{��1��#���UC��z,ԌZ�h��.z�Th�8x�Çr]��uY�
����;"cZűtn�j d�-x<�K��ӡ� R"ό�=�J[r	�e�Gh�$xۍ7A�V��iNYK�a2Xۄ�>�7m��춱۳��j���o�|���"� ������!��X�����PzR7&x
�,��p	/�Vz~F Xl"��kA��^�	;�<Z�?.e,�����p��'H���t�-��/w�b�� ���աk�đ�*�	�}����o-Eg�+J��K�w��s���31�j	@i��SQM0�^ZÏ봘^� I�l�a��]E9���gO���F�����,P�b�j��Û�䬴��8�s�A��� ��c���1�������,z3�;�2ϲ:�����ܡ���n@��lC��nX�a����'�:4��X6!�;�j�-ۛK��[��$3�rʐ��[����ۻ-�,fBgA��P�S�#���KN�A!���4Z������֖a�B?��ʛw;+w��x�'>�\�,��e ��L���2��Q��
Р:�A�z�C�����^
;q��F!���ՐF�Kf2��'�h�D���%��ǛO;�%XW!"I��s3�V#/��CƟA�D+��3����[���t��[Q3��"����Dyv'3I��n���l�%��X�3�����m?�ظ�����)
W��{�����@��(��H�ɹ�"i���_�Xk{�.�&�L�3A<�g-�4u��9v�tk�Q��o�֠��-KMd�.�v�o���C[h�A��H���[F���w�+���Ƭ� �귓,�0��T�����q^��%�b>�XtMc#]�%oN���S�{�-�T������l�<���+��ȏ��Z�@; �J������D��2e	S�.�8C��g4.�_XXV�b�c7�\���SQ�|��B�
T*<��d�)bZK�����U�m#�(�֭ƺ��]�*ڤaq��@�bb���1��E8N#�{z�˦�_X���y=ag4�4d��]��*�)|�e�o��6ѭ�	xHD�;�c2s���ݬ��y����,�6�����Q��x���\�?B��0f�_�S�r�|��>�sS�A��u���r[�����)�p׹�r8\c����(rH�����WA�9&	I@��p�;�󎇫K�XL�����j�oܓ�_��|�9b��'���B���;��8�\���q�80�6��\@~ �Kf�#Z1M�y�&3��T]o�#
b,��Xfy�G�JM#<��㫫��##��\2}]w��A hje-]+٤�gQ���	`�H��+!����mNHJg4��C!�^��Kl���'~ݴ��&ݢ3���x�"����ْz1����Q�>'
O5]���g�N2aȫ�蔘�r#�5fe��߬�p|;���zjE��pW����V���BW�3>�3}�����^�|�jmk K�w��)O�����|,�{�\Tܴ��a-�[���E���W���EzB�����*��#dg|F_���*8"�lDj��L`�pg�>�L�HV �ɩw�΋&�2!Zt�v�6ଞg�������O6���[���~���R�/�j����,��{,��"E4��Έ%)���KtD���0�+k��SS�f����F���,"RW9a��6�ڦy�8�`)�в疕2��$i�C�b+���Ǌ�ُL�R�FH��	2-��P/9T�gw���dG�z�w� �K�´"ּ�&��9&�mk	�T!�Qa/D*��D��!%_���{�u��G��V��]��{���vV�W�1��R�0〄(�81�sӮ�H�
��,�]'������	C��Lq��?p�dM�,�!G�>7:��U+fBW*���c�l
ϳ���ć�t�Di��0�4�6t&�NS"���`�E8����j9�U��>n�k����Vo��)KC�Ta�J���rg�Se��ٴ��ܠ�	�}��E	�2������@�D�\e�f����+��ݾ���DN}�j��MX��Ql�s5�:���in���#�w[�7�O�틛`Wj��������̀��x��6t�C�?�&�BC#X32�
)i�Y���n�v����$I�jO/�G�ֿ*�>�	 ��F˯�9��L�MC/��n�t���&_�|}���O2-/pM;8��F%��T������Dx� �[�}oM��5r�~Y�B�j5&��N7.z�ے�yY���և�uxg��4!F�_���eC8'�Y֝Dн㓣�`z�?�6�P�Ⴐ�e�]��2+oZb9���j�g�t�B���故'$�{�4�S��+[�;����k��M�r!9Ϗ�U�Lv��k�����7��4� DC�#�#����baUM3���U��
՟����4M��Z���[1���7���I�g6Zb�Ol�BI�&�`ln |�� H2��*VAmZY�)گ��T�4H���Aԏ�ۡ�E�=^D�%3wJ5�D�g�thJ�n�V�dX�lɈ�z�_G�Ľ6o��T�D.o�r*mz�Ms��
{�3ֵ������ຖ�f[�m�A�'�ǃـ�I�_���K3�
�A� )���dO?6�1���g�8���0���%�����<(���p־�bʟ�
��ć�����6 RR7���}Z�'��4u������yl�q��{��h�����9��a���9��fyՀ�Y`H��U��܅aa?=0hN=\

0�Dӟ�����{<>
���艤� c���-m
I<�qrr���`H�Í���8_�L��� ����#�=�rk�"9�$<T=t۞���8��-<�Q�\�j��SIə�����K�o?�B�{�b��$³v"�Kc,�蛷O�Dk�M]v�:���,��Y�J�`k�g0�M�y����	��/!.\��2��'Fo��j���&�밄�Z��S�u����)a5�cwR��ˋ<s�Ӆ��"��!�2ř"~�(٢R��:t[�VB��c�ȫ�Ζξ��_(C��u-���p?��J��4[�h�������
�&���ӱ?Mngx�P�㖌k��s�����>�T<��R�Y����2z��ՆZ�YcJ�+�L���̍��w|�!�nC��L-�^��1-�$�(��!~IJ���;�5���;]cMC�g(>[�n��힝f��b	\Q)ؖ\�=j�L��(R��$E��8�=�s�=R�����	��Ji�� ����vuD��܁�oo+f�ͦ��a�~ԵZ���e�o�}T��*�6�/iC�'Z�㔳�!�:y[�Ę~sS#-��D\(\�?��^�\������z���$2���u#bG���#ұ��o��t���g^��}Ɛ��K���؀4�	�H}��d�iX�\gm��w6�t�vpQ��.F��hV{-%V�Pt�Tj|6�w�à�T_*F0MN�W鑃�L��|&~ӟe��(��/���h�{��}:e�kJ�>p!�jȺ��O{9[i6 ��M�.���M��W����(	x�j�}��p���>v����.w�m�����-<�u�����@�.s�~L�}�K��0QH"�]��ΥA }�f�6{��7S�p{�K@��2f��W¤P���g&#���ׂ��퟇Ӂ�‰ku;fy-�Ҧ��������Ց,=����5��3�Y�S����Ǿ�+_�3�z�����
?�� �$wH�B�~Y�K��\0PQ��؟��,>k��f=4q<�Sv��Q��46��e��ijFa�Z�xG<�Y�Q�|����^F�����i�C���~�a���c}l�'	��O��%�Ƶ��1�ҦQg�	�--m床,Xr�Y��u�EY;��pc��א��5Y9�_�ڊ�)f�[�[�%��HC��@�ᢿ���)��P���ʠ�V����]�;�� �FW7�bw3<O�qi)'���aBi����{w�8	�p�F�����Յ[;�bA!׉Uv�7�s�w��dQ2��]��EM!��]��L4������X-���f 됻Ke,��� c^r�<�#�V�i�/gf,���Oy�$�NH���gގ��g:�8�" �Ab��E Z���Dλ
��C���ti���lu�?;,���XY|�����.�c��������%�(��w�d۪אw�=�;+G�W���d�NC�AvQ`\���f���ޒ�򹳨�l�M3�4:�kg�D;�{����+�L8+���K7�g�a���=��5a��;��=�ӟ~$ֽw7�e��al��x�ā��Z�Հ��Q�29R��^�UwjNG��HC�~��e+8��{���
����*Ee�z�a�t��|�ts�U�I�(<f��~�P��i��y0��-iަ����ɁŠ���]�B��F�DP�kl�����vݽ�5�]�N���Cx	}Y��#ro1��\n��r�wP{R�<x���� h�F���b����gOx�����Öٍ ��j���
���W�j�J� �<���m7�I���J��)\�2Q6"S�I���W�"·^_8�f�������F����SyK��U�~Yw�ACG�8�$��8)��9���ɪ.��ae�s��"��3%�����H��8�������4�Wh|u�bq�3%���.���lnl�"ƌ�'���(�K�	�n���)��B�N׊���7<���%�P��t(h#3ZX� �?`��|l�trk�Jx���)��ItL~��eA!������=���RT�ɳ�z%�E�Ps��)�u���%�9���!��ڮaKK��b�w�[@�$p�Gj�HB�2�����>O�������gu��D��kqm~���0�̨P����$��R)��9Xri����3��PC.F�6%�1�̕����� ˹���E�� |�A����� ���	�|����,�#:B�~ա���J���E�Z��Z��41�D�a1���]R!w��sf��I�*n�ɰ��q��z.G驼
_>~�z+V�����{A'�9>jC�Smy�x�)�h���M�H'�C�؇��Q��F�=��A>����Â?�*�9p���e2Nw��'WQ����:I����K\��E�++4B��'���Lt�������j^���a\ �#��
ˋެ�J��a��-8�rrx_ĠA�Ma�>��wc�����t�4Z� /֯$nl���w'rQ\�b����ѕDbrej��̅t/L+o�����y��t�%����n�a�����>I���C����ݗ�n���z������^3Er~m���������g�v�=�RxF#30���9�w���j�f�"��Y�_X�(n�XW1g�K"C����W�T�Dh�8���槰�M�F������2�2�H��¢;ouD(ؓ����"�tMC�z�)�xӌ�,t��� }��{�q�:aF��b�R,�zD�pђ5�i���"��b������ĭ0�=��yb	�-����@�̒�@+�������M�Q<0�C��0�T�7j����k��0fG��4��j߉b��h�Gp7<p�c;�����N\�qbx6�����h��I<k�M����4��0�G%5g�Tv��,��S�ؐm>-=b֎DTg������\q?�x�h����?���� �����7������f"xM7,&�ϏnvMʙR�=81��8�����z��^A�!/��c�Q�z����,1뤗��[�L+C�qM�@�)��.�7x���2��1���I�o,&�W��:�8bI���礠�m��LO�:k�FD�~�뎢�{=�;4a�L�L�����'Z��"1P�9CN�d�6�a���O�{x���xA�9�a(�M�g�������o��{f�q�G�n�F}~��*/�,RS5���̲x|Ғ�rV�)�z�XӐ3T����g��T^E��M�(���5����W��[A�d�/��K�4W]���&����p�f޶����F�Ĝ�{^}��f�S���c􁳔�����w���~����4��X�]��|q�a�K2+�}��G ����xp��k�D��������p]��.�����R�G@W��O�Q칣2kP�v�pr}����9�w,%��.�i#ȽeC�o���Iy#zD"LԌ&-�$�գ�s�{��W~<�M��L�m���\)���ێ�I��瑂����`�&�ɇ"�8�7�ڣ���}�1��?�l����Z���ҫE�mP!X�g�q�����^�ho�J!|Cĭ�(���܍�W1,�$aV=�m�&�-���nBN����D�e�\���N�r�*Nv��?8o�fչ]���UA8F�e1aA_�Z�z��ً~L�c��)�#���H��z$�-������L���_(|��E��G'��/�������D#���
>�23��{�R'���W*	J5�N��n곃h��qC��aMn���-�9ς��:�.k���E}�+�`�W5n@�����E<��KŹye���9��l�)�����t�4�͌�V3�$�fL�黇V�GS9;u�����w/��F'�t�h�]L����ly�����o饤­�]߳y,�ߘo�N"eeI���l��T��d�v���t�Gר-��WF��b��vM�o��`t�}�s��	-�gNhIό��{a#Q��kK!��A�v��N�sy݁e�5���c_�`6|�P]���Ʉ�	|~ �V���4������+D�8�Wk��<
�:����� �ӌ��I�%F�2t?@�'2fq�E>UՍ�8j���t0s(�6_�J���i�J�d��;ZQgˮө�h����tw�A:��MG�ӹ)I�j@n�&s�f�	��sUU����2�إ!P�h�'O�s����W��f�rZ�hu�0`���V�H�(�������(j��!>�7'!DY��Z���X9�2 �m��j�AR�!Sy!�Њ E�Z�mhb#��xd����R��Y��/km��g�/���x��ܜ6�̃��6�H-�UU	��u�3���Rg�s��Ґ�d|�8T���C�o���-誹��j��p��yޜ+P�6k}z}��x�l��[=���u��׫P,��O����5/��bH��o�n"cԥ�C�E�W`I�n�\����G�+�%8���&�]��a����[���zͅ�hh	���:���B���.貌k� ��qsr}Q��Z(|x/z��n�>��G���}�n��	:���߀�n�p��{��N��U���2�G��oM� 3-33|��o{[D��KM�����&��s�^P@x�OpH�<�#׀�X\U��L����t����Ӄ)��8H4j�R�6%ph��	��i��$�K@�4�Y.�O,f�^����]gVUuo���j�OQ�m
oE��I wԣ�	��J54�BӲ?"|������"QQZ{�#�a�E]���5�\�
���o��c
W=%z F;~��)�s?�H�P��!q휉�{��Es�%i���"���
<㫂�#d��%���=p�u&B�-�h���Ɍ��q~M�,q,^~e$!����d��]�~l�+���Ȑ�ova�u��3��7䫄�7?�~��a-Z:�-:>z>���H�.�h��*;��t�pPgװx3Ng��m�9iO?� ������
��3�6�C����We��X��`�/�_PQ���jE-x��nձvJپ�@���)7�O&�Q,�ה�U69�|�Pn�w�����?=�&���9��Q��<�~:eRR�F���ǳi�k�>}��j=E1�ݝ�B��:>�L%�-��D@}�����H�T�4h��ʵ���O�Jl��bs�Fkܐceݥg�2h��Km�9+�s�Be>�8�z�I�ĺ�)�0E�?�'+f4����V�Iv�K��^����ę��A���Et��6$�Y��^_�uu�T4�	o�+󈞦Ʊ	� 8>J�21#P悑�1̈L3���~���|��^��)߆��%���t(����M,|��^TI�e�? :��UԈKb��[����tB�R:coO#�6�����O<D��/�\��ŭz���7%��51d��5�ޫo=�����,y�����YN̯�[{~*�������JMF	��<�<5i���,,�KN�( �O�ۈ0R�W%L[�D'�Ί�����myA���~R9����8m�R�~�m�G眕͜ڈ�p:�hc��u�=�9@O44�c����K#M2'K��F�ٚ8D�\
Ң7�?�G�d�W֝%�ь!�L�	��������<ϳ^�2g��t�y�
�����$����'��'��4���!��1>�b"C���`�,|��zJ/53��ڣ�K��<���.9�h����K����.�8u'�vۦ�3Ӻ�Ҹ�F���g4Q�XK�u�be��؈퇼�����H��`]�[ae�D �xv�q�S�h!�!n��)�y��ђg2��{�?;m��ǂ�1���
��*�6�����-꭭�{��&�����s�z��b��B򊇯�U���	sN�)�sbռ��������uo�Z�dR?�T�6�%S::T��\�B=3�GQ"��/�ٖ��� $�rޟJb�N����j6��=S�Yp�ugY�r�2�	5U�"g٩	�w�̀��\��+x|�	���N<������ :��_�0�	����-y~��u=�3,��QR�կ��m�>�3����4>/���@�5-ؕ�^�L%�t~C�N�o�Q�&C�3l���R��R�U0[j/�H#�;����Q�-?�vD>z�╹���x�o�\d�N!M})g��s$Wy=�]+�FN���e�7�(]'��w-ߩ�ą�G����m([rk0dP�f$Kfw8@r�(0(��x/��+�/�
̍<&�ُ P^�2�Q&���9ER�Y7�h��6w1e��I���0�ФP⺮�5ˤ��d=x`�(r<�(��V��T�ś��݌;8���V���c8_���J ���E�9;��� �ΥB�����-�ؽb��NW���fYq߰��S�K���$�BXQқYN_4�=m��HYZ>z]�(�l7���+�f�(b�[��|h�C[�Y�����l3="�=m�v�9���댃	�\���	`�׷�Z��|N����i��1�������������y��Ç��J/C�I����� �r��P�2��@��KS��8E�zzCZ���v6��� �Db������p�yu�<�>X�uJtrǔf理Ce'����8����O�D�o���՛Xv��L���&��ށ��bs�����䳏�TE #��dQu��̮ٕ�*JzX�,%����*J�ߍ���ʄ�"J�)��E��8'��`&��<c�ͧ$��7���ϯ�\�wt3�],\�Ŝ����^��w�zrHlʔ��y�uF��'��!q���@Hv���]r��P��r���5�.���݆Z��I �0���&K�Qb���M��$�<����[�eh�ˆ��|��ʁ�e�p[Af��%��_P�m/�����AJ�_
nŁf�Hz���G�Dv/� �+�N<�@ڼ<T�ӥ��:h�c`(3�Nz����?��[��*֣&hv�h�Ȏ09�����s *�M�Rq�dN�����CϠ�ϵ)�E��٩��S1�Xу�]�x��,.�=h�<{�Jb%�=��2|L�u��O�����HM��7�]Ud�i�(��CH�+�M,a�7Z��A�s�tx2!��~�3�X�{/��&�[����j��xh�: j�vB1��f�����	��������,ϯ�m��\>`��<�#Ȯ{R)D�ns��d�Ӏk�Ϥ&��u�]xbDN��f0���J��9,������Ĝ:>���ȷ�|U�]�ߠ��	�I
N25�~�cb���u�v��j7u����JI���0�����c{ ��3oɻ����ߋ�kv)�!���v�O�ơ}�)�(�����p��Db��+Ռ�`}�6��^tDe��5��8�_�{_5��A�O�i�Q��G��T��H����'��U�0K ��PL�8��,�6�|�4W��%3U�:�$��[	�'�%�ۦps&H+A�%\9�]y�,R�+�m�{��B�Q? ��Ry�^�8���	��N~c��u�Ywک
%>bN�-W����U1J��n�z�x��A�8�{y���_�-��=T ?�Bqw�{w`����C�'���A�gZinη��GuBF�@�p��HN�OE�W*�HPN��WQ_�o����_�W%��R%�����b�]�t���J}f|��1��p��@v'�<�og���0�m�7_��!a��$�ōCE9E,�#WiØH��"�J�5��)祜�Gf)d85��aK<���q���	�(Y|�鿡2c��Z����uE�q�&�$��h������^2��^g��Ce[`b@��px��h�Ľ�/�em[�ba*�a�	��j�gY�S��/^[�� `�רX��1-8_7t߲���$�aG�kc�խ�*�׺�y�e����P{*%y��ζ�:4h���M��36�g�!$C3��p���_���[�=N�oRm�⚫�	��]��?��_����E>,+�M�����Wp���M��������|���c=1��Ad��W�"NsC��ư������������jvg�lX}�J_ +��y1?�R%�;����	�'�"#<s+�b���[�O�qݖ�	H�e���J
����R��n̓2���#-E8n�߃T�L�`�*k��ߪ�qЕ��"V��ُ>���D�1�a��ӛ�����>���P���p�ż�IuB��`/�W���@w�@��=�M�F���a�����N�b��T;BRF/�9�[.��(+�g�A�&��@��]r}J��-J~{c��=��H���c��1Ru���<�Z�
���⒕ah�6�9���z���}�\��g�1���Lu#�,*��u�g�it����/5�ʹ�%9�����'K�ѝC�s�����e.�W@bD]�����L�d��1h��|���pnvW��`�z9Łˆ.4]v�~��F����B-9�n��XX�v���F~�&9,�p�V/e����;X��-r���*2�]>�F�&�

JQ��p�Rp4�#䵀�4J��/��PII�\�R�+*Tr0*l1Ӱ�1]�}�M�*B)eɥu���� Ky�N����&��}��E�^��ʤ�@~a/�I&��g���� �3�'�SNfx���B<�l�C�<N��Q?��YQ4��GVu_�Ǣ�%+��ఠ�r��(m�M���h����@��Ɔ(RCb1�8�bb�N�O�B ���f��C�5�?�k���/}��RP	�f���i�ԳAV�5�!bŖ�xHt�c��	�J��>���	T�S_��i�3�r��\��gS#;^������
n��{]w�n����|
˓`�R携S`/t�|D؆XSjP��W��=��	TNY�a�~�TCF~A�4��4�~,H�L`�_����"��(=Yq[�9�A��H<�#)���A/l$%�R�CBB+���$mN���캻�V�7T����2���U"ćr�Y�K��a�P'!��Sf���,�<���x����	�qKF�.uy�K� l��wg9�T��#�Y� �B����Ժ��.�]��%T��D�Q+}(9��4�!�2�h�DH����­�>���i�!"�//eN8�u~=���� ��@9AԪ ��} �8�J������Q�y��� �; �;��.����Ve'��T�"a�LW���t����$�8Q�^V<���O���&�_��L��)�M3�����h��pNuz�I��s2O�2o� :[꫐�3���p�7��#R��Ĕ7.}ff�XB�/����!��VeL@p�Y�y�4N��)�v��]Aj�z@"*�=��V_�3���Don��ꢨ�	-~/��~��3?�ww��/�ڍ���>���B��~�ߪ�8�ߔ�@�]秤�W�͆7~�q�×�1�`յIB�)�z\���� ��]2n���ך��1)���	8�b���P%���û��N��S��$�Y���U�\�3R�y��WA=-�&�g��r��Ф]l\=�Ƒ�vb�Gؠ����.M�v/���Yp�3䞻s�#	���x% �TBo�T��.F9\�p�L���4�V�H����9M�+��ҙ�:�jJp)�'�PG!�m�]�h�ѹ��}/o�r�F�~���05r����[H���>���WP_�'�m-�y������	P$��vI�[�!a�<s�CH��,�$oܬ���ţe�D�:�����*�[��7� z@A���)0P|�B4��*c]��6_V&ke5�L6|i~HT�3��W�^&�݆��ʚ����9
�pCm���z���o�V	s1���p�Y/��A�����1j�>��S�z�υ:Q���x}�:ItE+'����l�'/���0Y��N�@���}�� %��Gt-(���+\��VMد�i�&�u��zV�S�kΰ�!��i��$�gd�r�+�LJy/7���5�k�;�&zUF��>F=�W�	ߴO	Q�.P�)�>6�\l���uەEž�ު,��ڒ@);�~,d�����8���,��(Ȅ����<���ɫZ���|���� �ł�3_dAE%(-�I����ۚ$��~��;���+[��ynhx`K�p�`�D��N��rd�����羜0&�PAD��W� �B�҈Q���wl�	�h�[
ˮ�E"�/tC,�q� �3y�8��w��.���l��ez�Ns>��Br�T���p͜mǸ� �]��d�b��0�a`�=��\���d����+�����
���Y}��!�CG	P�HCZ�"'��y�8����x"��$u~s��s�������|�����Ǒ�d<�{�>RIq����5^<k��3��^wT�Z[RrT�%����K�*U-�WCC��p���9�>�f�u}9:h�3�ְ�'���ei�!'6n����� �T�)���E<��Aۯ��gǈ	2��kd�~�
�#٢g<*��Ŋm	?������ސT$�,�9���z���[m��L�P �������sW�a����5X(O��RD`��rՠ�D�J��(�Q3��o��b��}�V�l�������y��\Y8@��g�l�£6A��+HP��i��%ˣ�i�]��;'����d���+��� D�B
N�^�|�8'�Ӏ�e��FY고N���]�`5���-4Ξ}��/D1�+DĺԡB��3����v]Њ�y�B{��~�w#$�=9�Qv���DS!,������dK��1�uG�'PГ"�Zx���A���wA�Ao�C=�KhT�j� i�	�%�_�:hV�NW�!u�4(�x����2���v8��E���e:�xM�(^��H[�V�x�����;7x����X�w����)��y�!FL���&M�䊮�âڝ[��:�MVNq�L1!�4Xk�#7I[ݞ�j[j!����ǜ���ښ��x�(fZ�߮�`m��m�?��hҥ: ��1w[�Qi�eZ�:7��0/���1-pŸ�1 ���K&�Z�'C����i�v�Ƙ@���z^�5K�Ǡ��v/��N�)�I|hbT�ߥ툢Rm��
e�$�����]SV}��E� f�;�B�����B���
Y< ��~�'2��s6)M��X�7�9�.�Z��l��$Y5�pD)!U?�0̀,bY`�X}��4;Ed�7�5V�g�`�Q�!n��ڳ pn�}���#���^|�$�Y�ȣ�vVcM�e�{RYCt��$I����Y���#j�4��	'J���~�Ӷd(��
�-K	�n�&Y�q��⮣mi�!`�C� K|����P�9f��]��φ�L�{a��v����yF;���~~�7�����ܶsn����"q���qkFt����
eoߢ7~*���[�����T#E7^�'��jΑ^�ie���$G�/�K���y�ú/��θ�ZkZ�N�H�X�T��掟��)i��%(�����n����o��a /:�����g}ݎ0�}}��l�&zܢ��3����J�h_�"P٩�Y[
b����_N�(K�[n��M��[{5:2�/�,B���@�_��·3�C�SZf[�MZc�rƓ�^�������t"��/(�$&B�Kq�k+KVN���7�Q!SVe/G-{]�$���$�e0�<~�����>���8���Ƅ1^�H��2�|0��U�5C�u�5o���������1��]�5X1��6�3;mh��R��\k�9��!��r��S�<��A����yA�KS(��'6��ɴ��2�]�T�q�<?���of H� 1x�,ZE\�����!�!ډ���W�V��}������2"��<�������=d�Xd�b#�	ƠEذ�
x����\)n�kI�߉�:����]|���l��Ԩ�Y�O*e��}���ow	ׅ��!ve����^Ƚ\�4�]�.�,��HP>J�5)!�9q8�#�ٺ�P�n�4\��,��ea��^�~U���(V�8\�g�Ü(��Qo_@�;��'��H�k�(Yr��%
��RY���T4� �*ր����3Js0�LIS����� �_E��U4g�sE����:��<��A��˔�:>���Q�)�Ny��2���
Yi��ߜ&��Ү�:FO�����kυ��-�#�T�}����ҝ�Qm�A�!ni���Q8�{��9j����<{m���J��f�
�"Y.0 ���M+�t$ي2���+JBJ�;�c�n.�nوicM�o/����D.b�r��A�����p`ɴN_0b;�%�3��Q�����IY�l����1��9q�|	�b͎�0���)�Q�XT�.�N�Hǧ�w�R�s��y�'5���r����=������y)`Y�~�A�̗u���)��1�T�9�tx��y��D5�E u�]v����u�
��&6_H��%�P�]+*&�ޢ\u���з��kA�u���2�¬�n����Ԩ&�r3d�b�/ᙿL?��c�4K����z�a���Z�o��g��Z��� ��u≓Ѵ�I;�!^�zIc�9:��Il�ރ�ㇲ��יUw�l�8F���"�~��P�K��k�8�������bS��+z�Vkj���O}w�mS�q��G��f֭���{�.��'@��j��;#]��EZSҾT�O݄���$��P��G�#�O�T�H��l�hc�&�n[=�I��gC�i|y&��7/�XtI9a�$���&t$�Z�Y{�_=a|YT��R�l��ӧ��n����$R�or2!N�WGx'�e��{��Nb��| >��Y�j]&/u�u� q�,����(��}ѩ�15wV#�N|���l���ٮ���H1�e���i���T������Մ>�w0��s}�&gU���8�p�YCŪ����[>9b�i8g�cQ%�[�~u,������DOu��b��M(C%�N��)F�qt��a�H�×,�!&ԅ��r]��ZO��E�P%�C.��8�ǭפ��$[���@<
LܝBzqGy�{�5�D"ʫ���v������������^�F� �̀�Ƃ�̣[ݳ�1��_ïo԰f�y�
��ӽ�d� r�����J��^+������6��R���;"ٖ:U�Q�1���?%��˒ǡ���Bh|�Z�^��i|͐������սC�B�P� ��CH> �J�F�jF]�E�T�\sM%Tc�U�Y���bD
�>g.<>~�Xh(�N�Ι�?M���)A�������@��dhaڼ�(!���`v\��=�Q�g4Y��HJ����_������ƻ�s���Y4�
���� up��W���>��l��Ya$�nߏ�N��U٬3�ڇ��
�y�d�;� ��D��!���T��<��f�7������Gl�P�r@o��?:���#^�_��YLa�����5�_։�Ϝ�w�+#�iݯ��^z�JJe����\�B��>G8`��{l)�!)��
� �`� C}�4���f�q�Jn�:C�p���_����贜����^����4*��&󐡷I�V�	^wrU��j����0h�<~#����b��6V6[s�ūd��~K�g�t�+����W�	�T���yߺ�T	G��˅� � :�@E��݂��R[1��8w�[��ݿ�t�
Â��ޠ���(r�U��������>�V�K4,��z�uM$$�c��?+��/������d�X�kO���@(�WL0����+��E���mi���t2��'F���&�\̣ў���:fE'��R�?T�"�B�\v�u��2�N���Vj���󪽆�#~Cvk���0�(V����D���i<�(Z�VH���_HGg�E�r��C�9����7�J���FFT�/K3�n��;�$P��q����@bm%rtǌh��;��,I�@�ơ�r$y���@`q�d!r���Z�YW�Գo|�/zR!v�:�ӆF6��[�"��D�).�dB6.fO�5QH<K�n)1�RM/Qʔ�(K�9��u�1.�4���^-f���/I�9"R&����T���zW{�nC��N�38��l����;�aI_�}�b=��5~�y�{��������W'��A	����K���{{9<4�~	�&M��pA�< ��h� s�
�iV/�#������
�s� ��\bS��b>瀼vd+)ٳ������JBt
 �F�b�{[i	�dr,;�Y�<�0�j<��d�*<�S�����p�כ�Xٗ�C�C{Z�1�R�����;���,��t8�N���v��:����|�Rn�T�騆+R�����?_x����,�*(0c�O������[���_e�Q��� ;�$��u��1v��	��h�M�u�jR#�F\fO�5ۛ���W�@��'1
׍���h��j��~O �O�-؛�q7;ڂ���ۉ�JЋy��ƁzO����C�D7��/��jHa��g��>î����Y�j���mP*J\Z�I����񈎔 ��q��X�B��ĉ��4�u=��+,��/?� >��i�����s����I���>����<�8��cR������O�|z��FZ��+��Z�oB�aA4\������W6�)L@�eR�\��p����׺9)	�'Dw�6�=O7J��Ӛ���`��K�/�M�y{��y��I<�Z���X��b�k� ��jy��?s�"BN�� ٽ]:�|�Z�u�I�����塗�J4���^��8����fe��H�\��	L�#;�HԆ,�s.�D*�����A��� �}�(kGP����,3~O˅��ۺ�:8	^_�a�Tc�Nr��jBÏkM�W��^��"I5�JP��%�g���vT�<�) ������E�<vއnۑ��Ц�dL���\��� ;օ�QX���L�����ZҴ�}K8^�~��������0~s�3]~% HR��vF�Z�_�����1q���F0W���x`�����z6�k�b��?��A�'h��{ˡS����
?�Ͱ	NW�!��;M�ɖܕ����l�Y���1r��|��iA^i�jtr3`�\��]C@(�":$�Z�����0�e���%u��|_bN��z���
M[x��u�9����b���Fs��5SQ�
�g�.��G���a������u=�M1�'5=j��+m��G��C~j�"��$��wQ�6'��+Ɇh��!vx�-3�D���P�a���8��ݨʊKBqs� �{������J���"Vx��~��x��U<��Q&8M5���0SG>d}_[������8_*(e}�B���\�Y�%]���4ϑ�ʎ�20��æ� ~�����2�)�P������GuV�L.��ƘӍ l�(��gH�)�rH�ٌ]��Ht�P㜒c���Fz��?�t�T�#n��=�H���ܑ��M���d׮�M��'�Ջ�B��kW�n����8IChv
zط?��
`����m��7`���o�����Z}8x@�1��{�Z���v�i)��IG�;����DU^o�\���ZV�89�S>Au%��x����u;֬�����O������!@zn�����.2���D�V��˹R_���.�ݼ������l��2Y��/������F�8�{/��dy��D��5�<)ބy	���8��Ѱ��/��0��r��� ���{mfؒ���L�fD�����y��B�����݀�f�?��s�~���-Kb��@B�.��W���b��1�(&@5��Z
+���������D�.�> �3������)bp�q^=S��-��'?P��G���b6Us�~Nn�d���H&
J%��B`�&���ݮQ&wҮ��u4\���/�{�FU����|T���c��}�Z�jK�w��̭nG��Tys|�BoN6�4���)��e���8�I��X�+�)���,3������B��c:�x���r�-�j���6��:����c�{���k*�}%o�kNV{	�b�-�m|���OU�q�ċ'$�ɯס�~i�NSڪ����^g������xH�F���}�1J�����y,Tc5q���)����9�b�3I����A?�d5�����~f��Ko���R"N�����̬D������,����:3Ө�/�����?�򆪏�m��v�a��b3}��]a�8�;s���~�Y_Z�9g�l�GuKyX���V��Q��he��KϸW�0�����q/ YE�R-�ک5;ɹH��������z�C=��`/�� ��5@�o }P�ŒX�8�n��ܙo�YLS��v)&+lX�4	��/<��R�1���`YAE���>�>^I�V��<#�xZ:f�C����#�v!�0"�&W� m.��ȃ/�|�eƐ� ��J~+��n����.�!KWV ��C�L|���`�x%[E��`�_¾VSM�ӄvP�H ���E��G�l�sa*��ҿ���x�7/�G"���@��ٔ'�<wd�Zo-��Q�aHϳ(�0�,8��ʊ%+V�������VnO�$����U��ȡt�⛞�f�Y�j�˝o-x T���'W��#�2�����,�m�(/�aݨ��>����PT��]g� B ��6QD\훒��KAh��D?䁥&(�����@����(p���M9�^��=z��2��5�y�dš�0��}2���b���Oc����V�:�����Ҥ��e��%,5U8M����'|SMm� AB�bcz��A!�;'F�gkJ3�i��_� N��Ò_l�8Mh[����G�7h�O����R�C8�i>?���iЀϟ�e�V B����?*�x׶lj���C1{���.P�R����{	��[�f��6Ά��w;�ҮKS�$7�1˵���Z�j��Y����ܯ���&П�`Z�}S����6��\�RPΟ>^���-�V�̙N�D4��;UL�_�m>0E�v��/x%�΁��H�Q��%�m@`���@�P6�5�뭨��1�U� ��T2$�S���K�T�"H�DVFI|��]g&�y5U7$M��9�Lo���2�L�47�����`ݎ�~�B���@���oݼ��M_�':Qu�g9й�R��dcyR%�n�@DB��G�O ���_�ꢖrJ�(U ��#�Y���"6w���:lW�(��NrlJF�[�6]�[�m:k��JN�#95E���t$p�䝼��T�_d�T������F�D��vj�#Y�?!]+a�ܸ�L�ǎJjV��0���B1�v1}��|�l�A���W��uB�Q!�s���1��h��C���$�-9�UglD`}�Z"���������J_�����3�lCo��5d9�Ոf�V�E�@���ۍ�R(�>?g)�L`�A�U7XD맳}��I^�v;Y�1��� ��[P��`����4�A��;$'[��A�0h.��I���������0�j#�*���b����C�]�B��dB��d���������FN;5�RNW1@s��i��PAaE���źa?.5w�L��A*
x����8���$.y�����+ݽ�LC۔b�|9�PL��9"��.o
v#
��0L�#��|��f����d��S%B)s=Ӝ?���KM���%���&��S �= }^��<@6#9UJZ�ݱWB�n������j�Fq�7��#3��/1��,6|u�0U��%x|MDz���%n˿����r��4RIz�1]� �L�VrXҼ�6]�IV:�v4q�������س@�r�P������X�����ml��k� Ld�K?f���s||C�����)�);�^(l����F�\R������D�M�ͱ��_�:� ��p� �-ea�"�NN&ǀ;<�a�Gi�Q�#� (|nR\R9U���PVX�ͷ�V �l���a�M�n�˶� \�⣋���y�*�KPm�6����<H��}��
Mf��¢H	N����9
��GXog-:�g�s@v�\�.e=���c����?@�H�IF)Ú��G��F�U�'{�\�` ��O�J�i������`�8��l%;?76 1B���#���>wca��m&�N�y=c�gv�|=��Е�+o_G'z#��UY��=�d!���bJ��ຯ���S�YW�4��Q7к�l���u4Wa�v_S&�lLı���vM���D�>��Q�
���E�{K�M��x�yP SaK7r�U�+s�B PTf>Aux��T0ŋ	�Kݼ5X��g|� ���a�����p9� *sw�?��X���{��1� ���$9S�I���$�-WK���٥��g���Z����\�OF'�ܚ�Ӵ�wSA���4d�(&�s�%lIy��i�V�Gh1xf3X�2�� [�*�rm��i�����G����}�q-�
�[�.�F�=�wřj��|��z_��:JsK��T��I~�����m�/�ܮ��ᥓ"Pģh�U�pbz,��wiK�An}��s�y[9�B�Z�k��x��T��K���p!U��s�**X8��粧�ߘ;Jv��_O�sh�n*g���<3߲�TC�:�~+����z�D���YI���AT����\�lT����[�T��#ogDU4|���w~l%[�F�n���9C��m벫�x�[�!fz"�^�щ�����qt�[�)��[C���L�s掩(��ݝ����ݮ�3]ڴT(�h�+�RM�W��	-�V� �|]x:��Fcc{z2"j��o5�I׏ғ�r}����1qR]A�GbN-k�>�0p*�YIְ}'��u�&l��yT$<�ԇl^���}D�kT 1)�zx��]ʊ���܃�o�Jbq�4���4H��[�1��-[�d*WO����I婴��P~ɼu' <<#�X��d�_�u���$	�y��Ѕ=�@m���G~�������jMN�+��NF�����Oh��	���$��T�\��'��UM㎌�����O
W"��!�
�N���ZG�\K�Y����%}x�O�2�b���?��=�(2|V��0v�pa=�<˥	�x��j���o�yp����z:<���jsp�;E�	���Џv:-�����X���O	Q�s��0��k�w�o'�bJa8�;��8)�=�$?G"�d��&λ��'v���>,�I��b�7N��\��,��~��%Z���zN��Z�k�*Xnn>I�2��Gۘ�-L�C}�NӠ�	@w���bZUeũRP vT���b��wɟ�	np#����*1B�_����%��˴2/r��4�Q��J~Bk�Og���vV��茂��ən�a���'ɉMc7`u�U�����4��sk���dK���k�c�M��'Q���u�3i��6�@B��{�)FP8����+�.����d��Fm5�s���Z�k�wF�|���tn�vyI9�T�#G]��i h����gBXP������'��лv^k�������E���: ̠�5٘�yRj4��n38l���.�e�s��-�3�Pm�r���C��f�H_�	��X�&j3]4N3�^|F�H~�ɷ�1l��W���/��6qL�/(M�&��7�q�!JŐ�3��$��,%��������J�򳖓p�o�B��d0�.�:��^�pOq���ga���D�1��{9h7N�8��'ʮ����LWc���EddW����ʦ]g�枕QC�o��	Y㴝./�m���G`���D��Kt;+�0Ժ�����\6Cc�ϳр&w��p���8�b�H��*�<W�Q���:s��^�����aY�3D=�[�Z c2v��1���%W�pd��t?��V�b�*����Y"��1�9�D(�����r�*ۓ]�kh���I�#cj<rd��W�^^���*л<օi���ذ� �0i��rE{ݧ��Rv��Eo��[��~� �>>�@*�4r�t@*2�`
�>�A�:_<^>�����R��suj�\ы	 ��`��5$ %-�E��ͧ��ʜ��� $3�G�&(���R!��ӠÐmMsK�koX����U�Ӿ����&�Ma1���֧t���Սv�T�u2��D>+M�-��m��D������е/�d��c�&ud���dhyrcVY��'l�qi^H�ǫkkeDk� ��M�:��5�4��]���`�ЫV[}���l�)�ޞj��!�L�/�/j�Qr��nN��(+�4NB*��m|]J���� 	ڄ1���30�����':!����8��BM��"���Ic�L�j�-{�nt��8D�8�IT�<��
�LIj݂y���W�������,Ŧ���|�!�����}�׆�Ș��Q�{��r#��g'~	�q��\�؍���o��B�lLm);g~e#F~k� ���t�sM����f�]7C�-K.æ����3=�HFA� Y�\=�נQō��_�Xd�y�5$�͉~�k&��Y����_�0��Ͳ�����T�/C��iVJ��N�Z.9ڣ�Ѵ$j�o���rO��5mZ8�$����T���S��Ӌ�5
3QK��K� |S��'[۾����m7��H�V���b
�E�>&s�y��: ��69pa�^�Ŀ���kn�{Uf���ا�b��a��������.
��x��A�+��ylp����������N��9!�p�O5TW��L��m�O��/�+���`l�ki�� ��QI��c�?�}
S������M(�Y!�S0��Z{[�4���P���v9F�����Ƿq^8R�[>�^j��xf�QRBH
,I��L���ݦ�WoR�d�nب�,�ށ���D(�����v��{̄�DК��R��!�����͍:' ����2^�-�/���	��#�R$V��y�e�|&D�f{-�l���"�|Q�b����2�̧�8��n��n�ݗLl| \N�A:��n��ؾ�ۭ�%4���zb��0�ȼ
ю���m�H,O�*�y���\D�f|���%��y��D����'��wb��-�4t�p0��3=-�-s��'�ya�(H�d]�,�*��J��I��T@�|4�ܠ�姅WW�5����M��N-�*�@[M([�+~�5�K�����ݶ�v��_�ޢjx!�Ǣ��3�Tph[�����#����.���R��{s*�*��%�1��3��@D���.���-?�����B}m�w�\�y5��5�Az�rE2p\���� <f�>�K��zt�nx�=aю?'���uw��U��Z�=����J��职�R.m�Yˆ�wW�@�/�}d���0$Z��`�y�n���,��O�ĸ�~m�a=�E�X�B���+7�@�K��Ppe09g��D�G�tZH�~�Զ��DM��؍W[��wW��D���+)�`���3�1<;XMG��-�$�I�ݡS�b�M�� ��1���{?�ցcݑ��uBP�+GA&R���)��%-��\Q�$�c�/��6
|oe�l�1��^mu&ϝ@sw�ю�_�b>�Q+;���u�A����P�����"�i�*eckW�r�� Yfe�G�ݢe�J8/#�_l�a��[xiJ	� �	�r�o�e����{b9���3_?� �|�P�uT���o������g(bN���b�K�#u�z�إ!����`F�1V�d�kGN�K�a�sk�t�b�:�"�m���aR�Dl�����+yA�	-��B��9Kѱ�5t\ջ!J�靆˕�a��O��T�-<1�BQ�>��A��Ɨٳ bW�E"�tN�Q�4'��r�Z�փ����=�7�*�	� b!��x���;��B��Zs�ˈ�����>�
��� ,��R0ĠN�*Ŏ�7F��^$-U�J�m�_��A'c� 9��O��S[�F���;�:�g�ʀ,�?�V�X��&�/`@���]�4k`� RQ�c�`�2Jr�K�i�*ٻ�J�A�t���roZ]o��)2r��ɸhH���Y<@���N��L9�m�BBh_+�{��W�zE%Ĉ�?�ҭ��)��*?m���/�7U�������@�V¡6r�ĨY�E�X�EaOt�>�;�%�@m� *$Ԥ �k�dDT5���}��0E�?�^ܮs��8�y9BFq�㰢c����.؝"�<�&�w�i�6ck���Ң�K�{��0Dn|�p,_e�3P���.��0���� l�s�L����4j����'�":d< �����❂l� ��n���
�l��ph��R���M�� ������E���r�P�����6M��d�^_�I bW9�h7G��k��@D�/Ϻ,ÐM���Rl��S�W:��	/��J~[a3�3Tb���8_<�`ǚ���ڡ�_3[D�8Eם������)P�E&�o�АZ����ӝWꗚɸD�B_���D����l�%�6V�,�l\K�#��e�1Y�$U�E0 ��"����2(v��H�U�@:d&cr��AK�Қ�:����`�HȚ�^�����iN���7F�Y7�j�����#���";YU���!��(�}��9���t��3���c�\����C�����S��01y�<ꑒ�$V�
BʳK�BLP�}�/6j��3������
���3'�>-�@v�}4>~��j�wB���:���w(̿�����S��e�Y����=�7<�|���f��c[c"%�������������1��7���_�Ѣ7���aW^�W7)u��b7!���҈��V�����Hs0�����"�����CzA��-�����g�˛��y	�kB�r�[���T���S�у~��s-���"/��TG��#z�怏m�,t�NޅELO{��[��tm���ڳ+�\�( 3@�m��7�Fr6�PɈ���s�Nh�$Q�o�S>������d>,��ZW(�_<�2�U��ʘ)�!���1����W��TX
��}��9�a1s��y
h c���_�E�,1gl�tw-f�4�O��q�}�;ݩ����9S�����Y��oww��\:9�Hv`��_ai� @�\�3�%��cÛ��O
;K�f��ߟ�:bh���k=����W{!N0%圐�5GC���Z����5���Cr0ǋP���r�7��M��pn���UxC $J f`�ɺ���鵾.�<Zz;��_1u�Yg�(l�aW����{��2��ⷭ~`8=s���8�.�G�6��KRc���v�mؿ�P
��!�Č�o�ݲ"��!U��n='~8*�Ua �0�F�`j�ңY�}c���g'���Ҥ��!��Y������w��
� ���p�9��TZ�vF�ɺ��܀a�Due�9Ʌ���t*��r����.�G���S$<�x��K?���/)���c-Э*�ث�p�P�WȻŒ��e|��6�j��i>@��>4lI%�$Q�Ч��}w�5M兣D��,�
N�W��}���'$���l]_�IP7��"�*$�>��^;�F*'��]Rk����k��lfS��*X��k����x��Y�u3�S�^P�K-u��)��N��E��?y"� q� U*1�����%0�nq����J�Q�q���%�cu��9�2��7r�'����h�����߿�*t?�G����c��b0��zo������H�A�ܿĩ�t~�V�I��u�	��3�E�؛�9HUk-�`tԋ��B��Ļ�H+��� Zu�hY^s2���%�M�	䍈~�~���ţ�WQ��#��1md%��Y��
��1�j�  ��;�.��2���NP���H(,�:W��P
��h�%�����l/���B�h2�oY����-�w"��X~�^��+����y,��JW�}�f�1g�C�/�	�Ļvu��-H�/C�n��a���R_���@�L�������UEwI��o�d~�tb6z?$��0�51|���W�@+/��+��<�0t��qϗKN!=8��kZ�L���Nd��]=�n�����N*!o��p���
͠ވ�o���b�q�d� �hUD��n��S+�Xd ^�&\s��}儮����	#Y6�.��gF#����u�Y�}U�����ӥ͙���Ӕ��iF�f�n@.2���eK��ON���?���� 2'�x����u�ˁ�r�zϰ��l�
D�����C�܍)�h���y��C�)1r OI��x���D=(�1�����q��D�1K�,�|�9��ɚ/�˖ �f��6��C��9h=@�����u���8��&5�K1�IƇ%��>?A`u7 ݱ5�G�E��;-�hIc�����*8�	���r��[}����ee�xX��5�Ә��%�,�R��7��$��ɕmK��Ӭ��q�G������?h���F��(��f���m�/J�P�ps~+ ��̱>wL"���<���:'��pXVڑ�6�j�r3{�O��`��ڸW�'��4�k��]�d�q�^�K�d1M���q�m�<ma�È9F.���!JA1d�^6��q%P��h&\`��;>l���Q�A|Ae&��,�*�L6�h�|?��Ӟ�]=���o4�r�(�睩2��!/��	�� s��c�=:8��ߌ�?f�倒�{<�ߤ��gPLw�tD_^G�޵�A�i{�mw� |Q7�=Gy�@�����ڀ����|�M��7[�0>\�0>?䕘�V��R�U���i���0,���	B���&�L��U���
j5��'�9dW��7M�H#��NϢ�w;ۀnL7�hw��oIy.<,��$,�Ez�Q ��x�0z =�M�|��.~č���\'�H]x��|uл
dp����,�6�2g�g�~`�����jA�l%��:-t ʣ�SX��	۟������ؽ(�S��Ci������_i�f���m_ O��'��=9;���WFuB�."ߘ{9��0�:Jze�U,	��-����b��q}X����\y ��˨����[��C�۩�'ߛ8���S��Onw���3�s��:� 9��@��{|o�`B (7�{� ���D�M�,�������5��]���X-Ã*u*�=cA#��I2��N�A�����/i�k #x�a%�%��W��L>��Mq�7�4Ƨ��$�������+g�C�$��
��0T����yx�Ko�1��>hqso��G˝$	lP�.����T��Ԙ|��k<8�;�����=�tUE����JN���A-Yf�l����9T!�~l�&d�
>�����r
;%���lIz�ğ�:iF�3��Z_iv~G�����#q/�&gbvǚ ��UE?bGl��n�����?h�fG����wq��\�hx{k�剜��������
���%:�C�MG��}h�FD䠀��#)��g��3�om9Pa��ڑj3FR��>�5��v����}H0jJ`2*�+,�c_~gi���clO��������ѾE�竺<6B��|�[
���$�����sX0�����I���?��_�^���i�b�� 6rNO�![Ā��\�ݳ`\��ժ˷�ƣc��l&ݏẃ��vX�G�:M�Q��,��(��<��X@�X^KvQ�}�=y\Ɇ�*Z%��5L'�H�j�f4&��P�����NÙ+$��V�y�%o�]�����v�>IGK,B̠��g�a��S/yS�K~�ɭ� &)��Nظ���)�@�E�Ұ$V!��;7iS#��n�xx�PKM���# "I��
�s�h�����0Ŝ=�����o�����]�V帖��ư�h,N�{� ���}����3�cB�z�
uK�4��z@ D�I�̈)�[��ۇS&�e7�"u�xb�^�X���B�ї�r�H��U��w�t��9�=d�V5H�#�z�yBX��������D]u�W�R�O�����)�nA�e����!�v=G�=�3�w��<�9
����b#h��G�3�:�^����H�I���L�#B��Ҹ��ǻN���w��9����L�� L�+���uϲ4 t�g��Z���t9�;:�"�>^�� �5�ݑsJ�7�H�I&���}��p0Y��?���۞<�ׄ'/Ij?�f47����a�b���]���.^<|i��|�Zx�:=�,���I�Qx�%��c�3ו�ߡqϪ(�_���Q{�N�c�f�{pW�F�����B7�Y
&-��C���xT��Aa �ܒ!"�c��=/Y�W�x�=iǦ�|+8�j����s�� l}�W+J�哀�ws�E/7@�Ŧ`0j�.r��H�eGi�j��������;�2x0�|��k�����N�����઺u� r��PX<{���c��!l��D�����%�Kv���\�����}^�<���)���ڙP|1�ړ��_���P�?�߷\�7���e�H^ �ͳ�F�qM�:�Tso:;�c�ݱR�滛|q�����#�hD'�c��re>>ES�lqX���C�|G���p�`�Q~�/٧ �)ь��k3^!�������|���.�CY��C��w	�.ȑ��Ñ���T��|jA�?Ѡ@��ů��6H��v`N���b9x��WRL�)Y���w���ׯ �F��"�!P��������\$�����13���h�,;FH��~zd�@�m�Mf�eW�\`){.�ě���h�5���7g��@߿'�T���LXj@ք��S�9��=`y�,��hIe���%Ǹ��DY�.Pag����j���m��eq�
��.������^4��L��+��L컄�S:H1����wme֯� J|G��� �\���<<{~��L�k�qvXt��`����Ew���R��Zи�+�o0nf�qז���`�Kt.�O ���9#�{�R�[t\/��?e��{�	�@��5!_x�E�#6�!��;I>�#�b����M�A�j���������:.L�+B�E�cpzŸ�:	���A7T�3ra�}����t�X���t�����w#��J�L���L�"X=O��.�Q���P�2k@Iz,b��5}��1Ѡ�x 4������6=29\f3�S*>��	D�gΑDwZ�Xq�6Fh�;��M��	�^M�5Z��s �%��*�R�ת�5v��t{�믞���3GN�O]�m�;��G�}@��,)��m
��&5ZHSH?>����wE6���[m-�蚳QN��C\���;�V�a��P�����m���Y�g?GT��|��ʹ6'��L�W�N���*Y.[Ο�[��K8G�
�������2ܚ�m��[�<0�͝w�e¯��+8D�8�jc<g�ܖ�E��{�G��x�_I�s+A��>T�������M��T��+I�u���F�������T�������n��Δ��������Fm"*w7����u#J}�9V���f�̋�`;L��j��L�u�C*����Ez.��v�Pd��9��z��M�.�w�T>[�Q�F��8���T����?�6�\��QL��]����<�F-�T��d �����oL�B9�X�D ��N���W�C�"iY��>�{��:!����O+[.���VY��Cw���U��]�R_>����㽼U˥"�L��a��Q�>��@HܓP�I�eY�v��;TW P�m��R ��l��<�LTP�`eǚEEU;�����5��C�h��0�9�a�|���D��-�T:�Û$X�m��N���qA�T��yp0��������$5���`���;��"��K�2���V���[2'd��?
e˵�o�
4��r	��b]w]��� �c����s�]�U9���fm��c4®���H��Һ��}���";d����nM�:.I�&65�ɠ�k��X�=�3V�2:��j�	�`�瀅��%�n��v������i%6�q�iʢ�Im]b��"b^4�O�$k|�F�+�4�� �L�b�DT���#�.�:~=���Fv�56����!ʄNkU2��0�-nKN��H�iO��u_���S���8��:�`}�4�$��c8��$��4wRɈ�&Yt���"�uTE�#e��x9t6"y���{~�h�+�sE�_����뒜�I�~�p鲏K˩w�7<���~W�Oᨵ(K�Yr�����v7";+Fs��DKl�*_�OI⒛�<P��7�k8�"`A�*C	ĸ�hjC�i4<;�:��l��ż� U~V`Q	���7J���06�TR6��­{�0B��G����~Y
�s�k�K�!f	ո��w+ҥ��g0�P�i�)I]�M�a	,\Y�M��1l�R��[~����2d9��������~��p�kj�砹�1<�@�ɾ'êa��Ђ{9j�a�A�^ѥ�4Se$��+�b��L�cCP8y7ݙ� Ȅ�L!���|F�5{��	��j�2J�|��=c�����9U�����5@��G�79 �)�H]%�)l�V1Zp��)���)zl)��l/ՍS�"7��rpvCK-����ʧ���m�Y�-�ڍԆ�1u/�^��)��o(�(Z'&Q`�8�I%����y���/SѠ�c��8+��׈�e��@!�Ŋ8�i�cV
����U8�.����,R���]	a��	VH}o�;v��;�wK߱�W�C}�,����n`��ɕ1r�J�[pl��UC������!�Q�|�w����ڸ�˻���mo�����6�c�h��NU>`�![�3:"���{�YB�Gp��,�>`V�V�=as0����fԚ7�s,�ܦ��[�TɄSa8��^R��0��QΑM�i(������~J�=�P�+�qZ��+p�|��r�ז�!e)\��.�TF��*rҮt�&CG�d��Z����5��ȶ�*~�I�l��<�����U�*�-{�u��n.FV�Z��74IPY1�SΔ�~�_��o��UxQw*ȿ��-?0���/��~Q�}`�Z5��5��[�_��gv�&��w��H9]�	�3$w�c\�#/�o���'��Ĵ�W�/��?���e���J��1��T�SE�:�Z�����҂����}K���Yt�T�c]b���j�WpyF� �@J�>�M�!�L�C:3�D�+쐧�3Y�c�Z�������XM��8 �G�`;�(%�&;���ţ�Vw�q?�N2�K85��?�As��܏Q���j�c�:�a?��9�ja��u�:Q+���4�E����%boޛ���d��q��c�x���,Gy�>�[ϒu��,5���d.�h�K�����}0��r�Z�s��|]޽�e{0��K�38�x.
�Z��v>��Ɖ�M�`�:ra��eai��^9�%��<'6���j@��ŕ��� �@���
��l�oK�d8�5�S]�7��V�5�eY.�X���%��G$�*-�4�j���W?��_����K���D��_��������/7����]�H��H��%��Ob�u��6h1s��u�<�4�ٔu��U
<�d`ȸ�5_�?@+�:bE�e�M�b\�n���`�9�'^�̴��;f��	.�K����u�P���ԕ/b�1!V0d�����peƠ���'|\���i&�������;�@�zͷ⍗�y�?
%�㔑�	��f?G��1��dN*��w�Q2|"K9�g��yxJv��ǭT#��N!+��{�	�"�.��RP�������na�H:��"�-�,����#��r 0���10��2K�QԗORg$�J��;�����xM�ZD
5"��Xk�V1>=�'�f�Hc9���5��|u6Ct���:k�t���bL�<.�jK6A��1����|ki��;��S�=/Q�u�1лI��?hu�������Z�6<<����0:$x�k��� &d]���!�Aj{;:k2�0'�x�/������wq_�&0�Y<����Nv��3J�4�]�	���rB�Y[�'����u�͠,8��O��+��h&�2����-�E(N�)���Bi�u���8����i0����)QLVձ#/Ys�QP�B|�����p��cƢiâ]�w�-X�����4�� ��h��KJΗ�n�b��|,�:~�_�8_�H���}=KZJ>��0����Ҷ�����~-"L���"�C��So��ú��yE?"u�h���Ǟ=P��HN�G.��uSՈ�i�8R��<ӿ-0��F�o�\� `��aL��W�.,h�.��<.��E5}�6���N�喇k�����R�qO�C��s�9����;�m���`z{�1b =aa�u�]��;���9�������4,2JJ�o�h��cp[�Ia��ӭ�y�X���%
5!��>�L,3��%T~'��t�rٴg�I��+�F���<:́�S\����)$N���:�4��=�R�p��*�[�MV�6F�f�h܎t��`��M�����1���Xn���n�~r�_�*L' Nn!�>��5�jVL��o���{��������b�8n~�=񢬅U�6W-�ݞS[w���8R����B;-�lf�vp��e�zH���RxH�U��x|E���0��d�P4
-��v��y��:frhp�.5�C��	�i�G
~�óB��f�N|��	�%�ٵ�����xN�OV��"��3x���R�� ���3��
C$��b.r��qj�����э����I⸛[_q/�����o��V��7C�:$�1ؖ��Zr��$�Ώ�ՠ'Q�f�Is��\�Tn�u�<(�;�q����ܿ���E��Ö+V��l���& t�������VH��u,��+���s�	'e	~�~���v�AG��d�U]IC募�nb����C"��s_�$ᐾ�F"�K�7`zu��$=粦���;(�og/o+J��k@x���\9��,Wo������O�f��`�0j�d���<��S����?bjڛl�������ɐ-���ۣ�Iϊ����`���I��ðWቡ�Ì�EE��8�y�z������?C�Í�Z?,���_(X�j��2μ�y�O^���u��4XX�$'�@;�q9�Y���-4�7@��Z���W^w��G���/���mM6�a��F; ib$R��N�ݝ�t@٨s��Hye�������~-���N�{��ǜ����Jm���|d�3�>�T?��q~g�Ħ��+d��P�t�����#��)�*�ҕ@,�K��eD���W_΀����/��@��W4�!�/8�(��&�t�b/	� DB79`4��6@�#�I�I��
QL|f��=K+�擩R��9�}>�O��#<b<�v�b�2���ӄ�y����B��7�+��u��1���y?@U�C��*}k��q�Bv�mN���vkx�[���ƕ�6����F��9x-�-�	�͌3���9�JZ?��ѣ�U��I��9n���P	c�n]�~��� �g����i���r,y�{���T[��D�[���Ŏ�ҵҼ^N�u���xkNESA��,�Ԍ<E2��^��\4a���2�(�`���B�'�X�A�%b�e����0�@�~�^�'�����^�\�w1�bI�O!�ξp���D��n����\e�:n*���Mͤ�v_n6�~P����}%͛n5�Q���"$S���ϳ(FI���ƈ��3!�~��-��Ś��=](U>\�բuGɍ�i�f	B
k�΁Pр�_}�2fƗ�%��
o������Q���K��b*I?��L�2�ɒ�7�NA�NB�3�G��V
^k���;��iJ+&3�AF��5���3�К@�գXo*��,3[��M6*�����i��BYK<9rU���p��%�UQ�؀L�h�
�p�u�1g�����?J u��(���EPw�d�E�č`FB���
���;i���j�P%d�lՑ��j,��e�P�A7F�T���N:Yʇ��;Y��`��I���6�Ή�?.e�w�� ot�1�*�~G_*��r��Z���e̤a-x�J�C����E���28�>{���b�β!�����b��/V;�Y�o��'pkЫ�h<�.�N}�:F��={#����|�q�q��A-KH
��{�\F�~=>e�o8!"��Hvkʰ�>ge���u���V���������֨E�<k�Qb1���C�_q���}��X"��_�Z7#��,�Vs�\�?%9���y=o;��8�I^���/Ve�U̲��h��S��m�"tV^i+W���p_j�-���:�!'�G�/.üq���������%٢��[�)μ���xu��P����v��ƘBN㜢J�+�?�;�{��H#a؂n�ͦ�h��JL�v�{�A��!��"��"[~裸�Pg�)����ޒFA�7�e��Tn���Lz��%eO?|��|�/~}�cc�pSE`�$��q���C6��GR��(��.s����� ��Ĺp�L���'V�[#��JG�v�7P?�t�@J�p�@!��N�EI8��FZ�	SP���n?Ѵ�E$K�R�9�b$���(��`#��(�'�$��_�ir����nT0�t��=e���8���C�t5��T�����/2��yH��=|-(.�����Y�m��~m��v%���XWD���r�%�Ʋ�Yц/�uCw*嵨5�2�eNdr�F�V̢���5g�ǐ�Ȃ#��U�/E�2�l֑�v�!�@h�N�K��c�Qg��&N���v�/�$�i����G�O��@k�<��g`��e8�g닧�K��@Ʃ¹ժ�T	NS�D7�
G�V��3��ˍY;&����q�Kh	t��+��^d��W�J�~�$�����W�]��t[:������DZ��2g�ץ�%t�2�ڪ��
ܘ\���"��Ĕ7<�g ��V������ű�I��}!q���?�O����A�"��g$Sӂ�,����Q�X=-N�鬀��#�M��_�"�?�(V��?�g\�hA1i�M���*0�w�8b��W����Ǯ�0��q$�*+n(1[ά��z���/�#�N��]!���������A��������u&ԤQ
�-�f���$	��.��53��P�Uj;ǅ�[�ңJ������"r�/�kaz���dE���j�{P�0+�_�#n�k���_�>+�%�N8�5.�.�[�|3P�^�t��X�ã�0�ϔ(2E̽o�vl��\;�2o�1����P���j�I��.�B�h����R�Ñ�	!�ݛ%���z�!��#�L	
TN� ������(�iO�?|k��~�Q��T<�>�ٻ1̈ a+�o�m�G&�ŕ�,a�^e�3���\
Y��o��pQu�>j�5�~���R?���&�	Bۉ�'�\��������@e��#��?�=��|�h(���?��ʀ��F�mڬP����b��oY�iA����|S��0շv�e���� �IT'F��e~�`�ǆ~lR��,3:'4�9Ra���
�@���|��q������STO8������@����&��AD���c���?I��Ԩ�	P��scїҭ+�mW����텽��Յ���7XMA��T�cƱ�!OA2��hù9t9ՑG�1;3�� =Ō�8�×�s<����������G�t&��=|{%�)0�EF����㌷,�@&�_}�w��������?J����ŐԮg�#��*�uݫ�b���|�A�򙓠��P�3STk�����#�Qp*�El��@X_��ԋQ�3�GX�i��ٳ`�[�O��&q��W���՚mq�=Ӕ�A���b��Isᐐ%a��K��2�{B�O�-B���'�9KTĥ��x�r�������7g��� �U"CI��]����ǚ�������S%���#ZK�Z3ڟ�:�N�����t����O���@��w�B݃#���e�pl�[]�B#[�������X��S���s��/CΛ8^W�&87k�o� ��s�� yԄ��o���a�uE] ���Z���\#%.�7 �)=э'h?e�#Ӝ�q�-V�ɛ2+�2Oi��o�a�R0�_.1��˘8N��SήO�g0h�{����|�f��$Q8�=�����5s����x�djx���lm]����Pz9�g�ͽ����02��	f!)eT�=�^�s��t�С~����U#�� ��'t0+t@?�O�EC ��6���b�R�q��]oڴ6��%�ƹmKK|g�[dF��Zb��u�#X�4���^EB��[��^�mU��݊$og��f5�,D���Rx����p̋݊�|E)0I��	�h4Ɩ�-����a��nI�����iZ؎��.}��b�G<�l6�Y�G��v��u�禠��l��)+*-��/T�j�F����, �#��F����,lV�c`=D�N�/�Q.��2�p����At�A���})+L[F,r<l���S�E��+��+��?��q�jVg��{�"p��O�˹��E^���f�~�����Q�F��Iq�u`��Q����U�/��>���)�ǵ�*�K�C(ļ�c�f����(R<<e�`s3���i�
���w���A���P�����*�H)�x�����i���O|�l�O����y�eh=`I�Kr������d�Tf�E��'�Kx�
	AZ\�.��I��ϴ0r�w��6��E���&���⹉��}1�_?��ҷ���s˅�$@��4��smf�}Z�uh>�2<����)f���P
�p�)�1��I ��4Hѭ�Os�+�X��`g@��ڦ��M��z���X�k3��R�V���G#M����j~�D@��*�-��%$�~-&ì>X�!�tT�v]��qJ��`�}����dS�6��*L��ycՙF������w7����N�*O5b��� �S%F�>'�K�JY�#j��d�Ҝ�Ŀz��UI3�B�)o��{�O���Ȣ���.V �~E��h��7ZH����������O�֥6�'|��h6�B�Vw���ҁ$����8H
���/���`a�EԊ�jt��Ձ�iUlOW�w�^��|�ޱJ\K���4dP�%�H$r��M?,��^�nV�?U�\ڈe��q�
�������2c����N�s.���(��dx>�*�Z��њ��X\��dL���$A_�Ω�q�xi�2sdB���Ş<ζ\gμ��!F�u��� ���#b������~=����@�&�FNH�1M�VөY25���J&�����	HT�8n��Qb�z�J/�Ev��N�_�F
�48t?n	K��qJ̔�&N�am)x���Dz���/�P���6H��P���)CGF+��-���0vƉ���A��c�/B���tQ��N]��;�����@����Q|�TS�nL3AA�(�������~JQf�:��R��ScpT��H�ޜ��M�����T����]S�wTrN�%F�r�8ϩ�����;PIyl�&$���"�<`�Ă1쏾�KWii$��E�f�R.����������]K�Ϲ�p�W�e@7��O��g�c��S�����m��bb�A��=X�G�[H}G�b6���L�w<�1������tPu���j_������.�~�vm�7�l���s�ƒ�jpx��
oɸiE�a�z}�`����}�!����pͅ~f�S�
�@�^t��d�e}as:�V_�u�|�q�6��?�y�Y���'����e���� �}�2UU
ƀm�!�q
�۹Ҭ���:Қ+xF��`m�B|��Y�����|s�&��v�܎���$��;u�^W�ae.��q�M�B��|%�|��̑�7%<�������֩�=\S���&�t�C&[�Qb>C��!zU�5n�	�R&�k�d���$�K"Bd�5c�l��x	�+M��k$�R�̈�a�R��ߵ�.�JM�4�Mf�FN`}��(��N,�R�	f*#�I�Z��S��f��2�.���th�?��0�Ϛ���o��L��$�|R�f^�͌�kJ��û��*��P���y�@�d$���沶����\B� )E�#v/\)�[�c$f��i5������^EmP�x3�}�{�=H�kk�>6���S��-!Pg����͓�,�,ga�ۤ�	��"09�Y���P�;?�]���f�2�{`Ȕ^%�ii9�P�XȐ�1��r��r����O*\�^�q�G�?�3��g
n�V}I	F�'=�!����0�ʆ�ul��o�X�йT��Bк�r�"R��|Cb���`&ڽ�Q��ղ0
���%�Ѯ�k4L2����s3�NSQ�Ut {�5ISR�|)��R���tQ�ԑF�ln��l�e���=�[� Q��,����w|�ng�� p�EQ�P5J�>��,?�E�J�4�sum�����xΕ�d	��4�$�� �6�%����`v�)��鶨e��
s����� �r�H��hN�7�a4�;:��N�-�@c�D}"f{'U5���,�iw�7�Iƒ����W��!dX�]? ��N6j`�9U��J���U�4,���ea��9���30#9#�郆��J^Ɔ�b+T*�5���d@ֶm�h4�/�k��\��pSFNy�_�5g�ٙɑ�c�z����#����cD4�&�	}�O�P~KO,ZMm�ȱ��8۾�U)�TCҶg7�� }�ڤ�kV)�.e'�A�4��!�_pU �Bd|�/*�,b��]@�L�u0�n��X1q��g�t0����}j���/&�M�f��'6�����g5(�C�������:'�'3]��3^�Ё�P[��zh�ÿL;�X:�kЕ�� ���E�pRP�;+ �˔�9�X���NX	P����U�>5�"/��z�f���_������h�+k�g�  @���S�1e �pk�y�|ntֽ�P��»�3�=B8�=#W����I6��߇�Hk�<=q��ZU��&ݭ�bꡪa��cq��-ě�n�a=N>z}�#�Ԫ��˻ވ��qA=n�G���n�.�h��YOd;�|ʅ>��f�	�����'����ٚCoj<ºx��^��e���f�Тd���- e\-�A]V��+M�Upi�����vX'���l�r8�u�s���AҜ���g̨�]7��H]��� j8��D��s��S���b*����*.������c�H�"�	A��6)���c�Q�VgL�G�7al�~��x(�u�j�Bj��&#O7�
ҩW�x��9�k�?/��?�Q��ʸ ���zq��PF����Wcf������:D�r��7�,'+.�W<���݊�P���D������-�̸c��.F�[�M��b]sY�/}����+1ףaY���.?�I�]����Jt�����gZ��h���VB ��a��Hk۹#�%ybF��ꩅ���J��$�!�\�$F�q��^E��� D�˫oZ�|������X�p�#��c�8Ś��`b&�ÐC��!Bm�9t8���@�p�f�����tS�I�2��=\�BE��&�x��+�5��u���[ce�GZ��A��2;������-r�m�R;.�;�h�-U\�}0�9���+�v��ƽFJ��T1���J�2*R��!KX䋢X*�@ ��z<`��2�汫s`�����#���6c�؊�{��S���ծ��(�*�1��&�C����w���$ʸ�a�����w�:��r3c3�2x�F��j4�­�
�$��kC�p�|���XS�(��� h�ʁbI�p�p��E��+�[��SɈ93|�i�zUhof�MT��.&�G�f��t�]���]jm=Vz4|a��b��@��?�g|��m(�apHX�o��@̥�{�Ϝ=e/Ø/K��S �ԋ ���@��A��4�����Ӻ8�ٛrKA4TP��I��<L�3�!�9h�{�٨Gx��k�_uUY��<�FW�O
LaL^4e1�9�U5�z�LG.�ʶ �d���L�y���2i-���V�zz��bzŒ8����@��O���?^K���0<�9˽�ɷ˞�f1�r-((̢����;�	}��Q�<߻no�w��q�B#�vB➋��V�������Q�]��T[\�W`|K8�<|����������w_$1��N��g�@�+#����e$��I��x(xLq�`Os*7LezHc�D�,P�@ED3�jr�	7D�*�<�4�s<�
�����B�<�p嬴�;T��Q�1
5 YA�;ɊL��JB�~��G��EF�������O��]�aH�ME�N�H�p��S^f�D9��b��_@X� ���_�Ezn�Vߝ,q���ousv�y�pϪ�c�I	�5jd}��9���	Ew��Չ��5n?��)6p8�`�u��E����P���k1�2l�g�v=���o���j�Ͽ�g��8d2慑�F=f��Ih�����Ɓ)����C�傟PE�*37���؇Y��,����֕�13`8W�4i�Wҗ�=��(n�<�В~m,�ٳ�̫I�������Z3��;BK�%��Y������b�u��{�� #�Z���Al�K�~������xZ��jtx���`�+�@l5����8�aw���n�?�0 �r�\W�6I�`��:�҂��*�pݏuq�{�FK���Ml�%?��4��VH,�����D<�����@�C&T;�{>���MΈ$����m��F'~�s ��j>{��%���) `�4�;~чQ��c%��%�.�woJ��yB}��_dK�?��0Pc:��ܤF�ؕΌ<���ܹc����K���d�d�\��H��fu�+�Ƽ�zܿ���� �b�_߷�:%Sv�P�/b�^'��']���CIH�$g������Sy:M6��{LO�Q:J�d"o�i��v-G(�ƌ´ܶ�tL�r񙓈{�´�y*ng^O6%�x�ߡ��)"���f��f�!���X�o�ȎY $�b��J3Y|�)+ 6�Z�=���
���mEw\-��u=3*XSh����	a�2��^��|S���)}��;��-l��L�6m11���g�7I��:�T��A6�9�F}"ؐ�D�q�yр���+��k;-�3��$����.]�`^ ՠs$�b�S�w��~�w�1�˃��0���a�����L���ا67X��8y�8X�SKh�|�-ylОvi�ۅ����� X��&ǉ��A�	M�/5�Q~*3?��ݼ��D��j�Sh�S7����4�u�$�V2Ѵ"���:"�Q����u��#K׹���V���>�zx�~�-��`g���Qr]T�Y?�+_`�a�~Ѱi.לyud� ���nIw�A��Ar�n�}	q}�ᕳ�pR\42?5A��qB��-St	|ѕ����(�K�Ė(��A�*�)�o=���W�2r�x�*�s�ċ�BP���=�v����(��g��B��OC�q96a�~��\�H�&�[d^'iB=��"�?�v���N-��I+�����/"&̼ɕ�0��[���"2{ݩ�S���	���5�o�{)$`I-�~K�0�M���Bu;o�1I���uE�����ȡŅ��f�7�t���&KHm�N`����o/~����u�����\�R��5v�2d3,�gM��{�N�i��[+���0��N��N
'��NB7���;$T8���lަ��,P9��	]q��&_C�g�Z�'�4Aҡ�g����:AZ���"$
�wGj|�M��/se����%��6d�������Xk=�Z�Ü�?����r�y� �rW'"'��>Z�#7�L.W:����=�p~���ڽ����&ظ���V��(f�Y� ݔ�*�P���^F3Mj�>�9Fir�4;wQ�f���P�9q?x˓ ��u������Ɲ����ڣ�I8�c̄	q��>���r�l���޾�� &�
W(�����W0�A'"~�1!��&Y���@��������!��ˁ|������&�pu�u�D���ñcs���w\��\�9�G�E,b3�#�UjO��#����~�XB��Yģ��S����W�rH������FS�5�hoQH�QPs�R������Iq:���%�s���7�5�V����>�H]d�*v�;�3	�H����n����0*�pـ�bQU�Uk�x�vǑ�F~y�Ҋ�6:h]��~CB����nj:�uhX��e'*{[y9WzIH_����R�8g�^E�vu"�>�۷%�W�}��/E�C�B��O�j��Ұ:�t�ɘD��_�Ox��蹡���/���k;miA�#9�%�j]�e4ּޮ�#+H�ʃ$%��:���t�1n.�YR2e9�僌��E^M���FB�#����b����Q3g�T9e���Mz|���PQj#8�~��ˤ�M�ݡ��M,:��"m�z�a��&XQ�E
���m-���)�Иk��ɗ<thyB2���1�*~�km���=[�P�nB�\�ɭ��;��*� #��q����E�����[�'fq9�A��~Nd!x'��ݩ]s>!Y�6���5�$�Z���;�XC8�?kP^���m�1��gtͷ����r# �t�Vu��}�ʇ�]�?�s�zwb���H������4 j�S�o�VU��#�?��F;Ċ�e�t��_u3/�
<����Y�8Jۘ:1���\�p�ڌ��7%B�6\�1�e��BL���g5� ��u��nr�*J*���r��C�zȺj��4�k�?�I��wd>'V9�b�Ov �T~�D@���c����՛%�r��o���c���*�5����|�,�u��NHs_���]�*ǡ�#B�{�zެ�'�hةy�$����������.�?�� �-(E<�["�>B�k� �~�Z��p}$�;���6�F'?.֌t�e�_�C�����p�T�f��Gj�;��:�n������f)v'#.��Bfp�1O@G��lt���;q�kB�D���5���&Lt�-v�孎A����z��=Nvڸ���ڱ�����<�.�3%9�+ʐCr�s��9��	�5foʛUjR��q)�\q�[1��	�e𬭚 �L9�JTܭ�O�3ɰ;���kg�n>؋����_QXZ�Bt<R�S��>��:rkؒj�o_�ص����Oy�F��8��*�W�Uq]{#�B�i䌫m���p�JG�^P���Y!����Y�= �e�f���E��'i�0z�+C��,^q�p�qI����L7f踅U1���VPp��/$`~�/�{wpV����`����g���I�O��KL2C�᫱.U� X;��+î�����2(�0ƨ�$�uo�W�����ԟjr&��c�����%ce��JL�ビ]{`[�ȶ!�M�瀰t-)$��i/=�Y<�ב��>a�]������@�+
�,j*�Y�H��T^���R�;qH��3Bu��`�;߀&��i5x/A0�C�	��f ���{��-�����#c�n��A�����.��pS3��R�1����H�\��X0"�R��i�'�-M�p���P�a�Ez����+�-q$���z�ҍ
���5�����9W�[E�ﶀz�1#=N#�ĮݝT�I�B���Y�J�&�j^��k���>�!����裦��H�X:؈�`�AU�~3!��fAb@���<���U�t|���Fe?ט�q�< �C��^��%�?���r���V�Ww�:���cx�a�$#�=�P�=����9�ڊ�F{���[uÈv�;��G�<}_�J�)ő����ƒ�$Y~�!���_j�պ�ư埅�Si�4@��S���������a�Yʀ �7�)_�G��J�c�=7�/!/�$��$nn�y����C�Kn�z��ߣ��h),�re��;L�1w�`L���-7�܃S��r��_k�~;�� :�3�w�q�+%���0g ȁ�3,UF���ո'����SK9���տ$^=�S�w9,�L��g m"�Bd$�����
�n�QOx�-�f�	��h��7P��t��P�"Õ��
Ovh	��`�p '!ʸ�Zi1O\�V���a�`"���B�s�6�&���]!A� �05�I���ӗ�� �GidF�OUD��2��8��]C���؎.��a�-��/�aE��d�U��ה�ϲ�U�\z nyY�b��_�L���dS� �j��>L� �Ż|3qd,~/G�J\j���X�Up~�Uɘ:��.^̰iN�����}j��jn�Er���CT�<��ֱ�#�����_�L'��&u��lT,��5���_�$g�؈�[<� %ּ{3�����r�����TM����,w��P�jV1)Aa�3@�Sd(1���y]������8Ҭ-FW�e�K���H0ժ�m�蛵QݸMCF�r��q}{��ͣ�u=T]�� �A�O1K������YȦVM���"��������jwcL�=���%���B�Ȅw���fG����J��`�p�N���fbl��h�_������K�`�JoX�3����\��H�J�y�O!�+��3��6$]�����"��1�J����YUrӞq�pn1 rѫ��v׳9U�B���7�.��HM��
���A`ğK1'���h���$�'#lk�M�kHw�gɘU %Z���TՉM^ ϖ	+"���''�l����޸r�l�c\t�"�s�V�G�x�����>�X.��a�M�l��!�W*�m"*�U���٨������Pg%�_醷�]H7%5�Cg�1��Ǆ��9ޛ��&h�9�ǣ���L�
�`m-R�q�ko��Xq#����g���L�I\6�|~&�O�� ;z�j�{iMF�T��8������ ~]wm��)[c���;�?O�f���>>C%��?^8n�$Bw^�6�S�>Yd\��È@��gW�m�zŉ�;Z(��{X3%�y�.i�1+n�G0^��q��! �� �V%�x�c�/4��]���8���[~g�_�E��F3rN�F�%������{@[rL���J�%ҏ?x�>����3��{ �����{�Y����p���CBҴ�[mLF��)��ݿ��[)�@����a�q5��t
�0)���Ҵ��++F�c�����!ʄf/��l7��"msC�7��"����lٞ�f�*'4����Tbڏ#���o;��2��}���9��f����}��W݁��M��uD�XO9��AA�=4�k�S�p�)"�֯0z��5���9���`i�1�QgwVl�܎�66)"�w�|7�-[�
l�gC�n�-O�6�rL����GuA36�2���0��d$|t�g�خ�?�����`h�O�@� �(�C��S�p��Beekд�G;�<�oZ��#�n�~�Y�u a��n�tȉ*��)Qo%�|����-��oU������_K7�b�Ȉ�Bp�?/6-<����{a��v"���'�]p[�3��P�V}��T=y�U�y���^u�H�aLT�ϐ�A��[�Px���Ҋ%��jG�|��j)CL�wb����L�ӡF��L��Uzkct�[�L\�k
~Jm)����h��V��)�]��#��7��*&�K0q�mf���HO�#�����R=��^@2�.'ӓ�z	˕��`T�a����{E����w��ߩ��18G���x)���B	�`A��J&^h5`:��ؾeXɓ��3�qҁ�{� � ���>�}�<`�����8�4��(�L��a��0d���`�#tm��)~��)v��{4���'��4�LZJ����fEDJ��7�נ��%�,�2�� a��y�X��<�{T|�?:�k��^<�Z��(���˗�b�9�R"������͙^EV����J��-FP�Ff�Y��g�b��[p���'�7Ju�j}-<�6L_G}O���9�H��~�R�7Pu<[~�+]l¢崈�3�M�pO��o��(=�)�z�>�fa�Q�xI��cř�js���	l�b~1�,��h)�_�5�UW<2X�I��7$��7�?�
���Y3@*@P��b�ܭ뒏�����+�&���V��g]��E�?/�of.":�J��q�0�7l�=�Q��9k�՛w��D`��3%}k#> �� �F�?+g>���'��A=��&;�{,��\�FrUg@v	�$x.ݛ/�͉���2'E��tu?]��[��=�I���KJ�YE�a��4r��w��8��:�0;[���h�8�vp�Yu����$b�4%N�"7'.���K�b-|��re���uFE���0kL1��=� �-qc#�C8��[b�)~hv���-�g�Y�>�3����!��ʂu�� 4Q��Np�Y�~��6�.N�Z�PB�I�A��cE��YC��}��z��!>�]k'4��fzKIZۯꔖ;���1u�:{j�/��V&a K^��O,�|���OMpBr�S����-ӕJ��ƢR��/9�o�ro�C-[};VMzn�jUZ�c'�$Zv��Iͬ�~?��kR�Dx^�+��k�^���n�Iɸ��W�h �*��r5l��\CΗT�NV�-?��ʉU�J|�Z�Ŋ�7}VK���}��*-exq^���z��:�{hX�[��y��cGW���L��+\�y�sh�p��&����f�|?�v��_C��~?��yk��.ӕyy��ӧ�!��O�;��5�L�<и'٧��o%K�&CkS}����ȧ�b�`��$�0Mj�U�A�6E8�Q�.�+R�O�)#�l+%��@L���h�~x>*�c��V�8�\�QV͍�֯5!��u^�w��s})����	�~��{Z�%`+��tfn�X�q�`����I�|y[�e�El��yt�S����Y�%���h��}BǏ+[������TAZ�,�ųo���JҼ�.�{&�5�\��Lmi����E�̝�db�Yr�G��R쑞&P�)w/��,��^�]������������)ԧ�e��i�ףt��
���'s6N}%-)mφB���1Ō�CN�o�5�
X�)��C3dh
���eO`r`^����TpI*�\�k�ߘ��VT�(�?��O0�"d�cG�݁�@�Γ��H��tV\���;�[/�'|�u�%(�,����=.u�(�Þ���ufNw�5ZF����Zꡌ<��Gqkrc���׺~��_�,����rG���ۉA��w)i�G����4�H3��d� ��ER�Z X�Y�aG�� NdT�}C�J� ��.����WrͺɅ=.T�4w�B��G,��jY�}���4��$�[fYt�m�[:r8�����Or.;�@�6��z2P�^Cb>F��x�����>	[;<�S	������HZ߭r��z�N��2�e�t�RFÕj�ɷ��?�EC��]�xQ�4Y�$�i�sc��f;P�A�+���S|��"�DϺ���h������{m�����B����{�@憸� aKQ
� "�,7,�!��a�d�WI��4��e2�ţ*��Z��x�>���/���)|�]Ki��0���4��$F:���;<K�2@��H��EUH�)�T��5̤�'�_��ޔՋT1X$�_WW���*2jL.PL�`A=�A`��
ʢmHSE��FF�����IpK�ӑ1s%Ef���ګ�h�W7c��ґ�}��\���þ�u�վ|���X�g}ԮK'+i��!]�]Q�u�$ɂ�\Mꋟ�s��j��"$'����>œ�4P��/K��=o�� ;0�R��?�?�2�W&�r���1%�6�yF�/�ϼa�4�U�uz^��<��`]��P=�.ut���`}�?�9���\�8�Z����H��,�W8b5�#�!�(w�����A�E{����/W(#h�����5�f纼N�GN�����/�۷�+d�T�X&����,����EƴߵO?~]���?����~��`�1�o���3��	��$��F�����(�:C���%����E[S�c!�S�� ���z�&HH���*�:XC�ZRW�A��t�Pb9�W��FN #���%f��f���Nߌ�D��� M\��m<��N�l[��^�&"���O��C%�XD�"!.�`&����7���xɢ�]	�b�����ō����΃B_����g}����M��߱�����@t,�C��{���~ԅ��7L·�_��N��=-
;>�|�����䵒��w��3w�v�% ��c6i7m\�l���&���J�ځ@�	2#��M $΅��A�?Z%����i���|�fㄋ�?��J����̍/^K5*0O|�Z�Y=�qq��,Rt!�1��a҇^u�Kʜ��G�<��g��ȶ���^*���+N{�~!]�
(ʠaP,�f���PꙪ����i/֥��e�m����Z��^��"������>+��O��g8;v�)W����y49x�+]�
wAU{��HW<��֘|_���4d]DQ)ZO��\YS�c0/�環��1����b�g��/*J��zR?�mdS���#?�d�>U�-E~�[tJ�9��N�V���,1?�Sc��35�ND���i���	а�@����0V�2������<Ϝu�KiY���M��4��������p�Zc�M)��_��ΙB)�K�/��Fihk-�����|<bc�v�,=���F�l9�j�MH5�Z����=|*>h�! ��6��ǀ�[�q��Z�'��l�e3v�1Jн������1�H1ľ�~����M�qvA��@��z�_~�����Y���cH�Ӓ[M����VѰx�En)`��;��:�z�L����SF�~�����2֐�� �d|�Җ����a@y5����8�3��[tϽYE%�;"�����"vX�-^�~�"�*QX���`��mpP���#���2-��_�y�f ��v��*E���"��R��b^k��tWp?~���Lo��L@�eQ��XӸ���@է=��/{��CW�z�&,���@?=���2��Bc|@���W�B�'$���n��eN��u�$��;;�j������=�� ��%����\Um��Z�ث��H��*o�����~3�(#Hut[�2�Qb75�!��!W>����(��ۓ^*m0��ڄ���+���7���%~Q��8�@p'��]��xT��ԗ1ˑ���ߞ���`�M���u���X���4����|����os����m��Ά�o�⇮����)-b�"�Ջm����tG���>?�D&.��,����S���G���hr�I�������KE𰙦J�X2BL�1}�!7DQ�GE
k�v����:����k}��9��(A���I�����1��ԍN��B�Q`��d��4!N_�G/���{�	�@/}}��K���؜i׊�"�Z���@�(Z@���"{��V�f&�6���ѓf�r�� �K�Y���M�xE n�f��@KzF��a}w|DZ.F�~����g̴���2��:n	>C"rS�u��~^,�)�aX!+8Q��7K��hӧ
���Jw�_�i�o?�,�n���`�-�Odh�Ϟ�¥'!�!E��*�x����I�@�/@ܥ�䧂0����Xr�yn��c]�o���%�Y!�%�[O��@��}��������_S���0-Pk��6�z��
�l|�#!�;y ���a�&�̦�u�� ��E���&p�-K�w�lT����.��n;����+LY@E)�Ã�?�,����4T1}�8��-&��(tيV�j������B�T8 E��Vg��W��	�X�����Or�����j �2� ߦG���\��#C'#�q5�� ;����$�U�T�s��`�s�X���ó��-��Ҿ�/JH�g���o�����,�?�Z��F�,�%
�L�eOr��Fߥ��8P�=}"�q�}��^�x�@���t�0���Y�|/ {�e_�lu��kE�E�.�D��p|����fP�����R�SO�����=�V��|Rj>�h�$�cG�׆�Q�a|yp�s��o�5��J�5^���B�ͯ8#��tH��{H{:��z��E��&�@	8/��=.��>w�z��/w}�kp��>�4[�_���'�&�:�)�ߥ���4M�+%1�R��c��N��(n"Έ�4a�� Vv����RT3%���*~�52��s30��v�NMW��'ϔ����4�tTL�QV�{t�o�n����������s��13�'�QB�X��E�ڢ%�F�!Z蔡 �K�>���6am��@�?�5�|�E8�1��[Sak���ťd�M�]��Zp�U��q]��!RѠ����� �I_%ֱ�$B�Z"eӏ�h9���)�OɌ4Z���Yۏ��X�M��sE�.�;v�y�qki`^��-�g6�nj�Z�H��Q�xP�����[�~�x�4E��{����.�O��n$����m���9q�T�w�*6����=v�x��L���@�k������E ��mѝ�����f�Z�Y[���Hn��{�̨��ZiA�2� s�+���j�QM�|i�l&���W0P믦!n�o,Ό���{���6���:��[��G~��L*��cY�?�:�sش�D��-�Ы��:�ߩ�����U�O@���\�F��JeF��]@ET���dhX'q�vG�^�g�l��베�%X�B��>�����+�a�3�2ʷ��&�.��4�2�]2]n���4�H\p�zE���F��X�Cvg��+p=5G��VU�S~d��1�R-vK#����WNi0�_ǋ��[��E���á�:mĎ	��̆0��Z ���8c�� ,��9%�mb�I\�uS���f�V]�4A���5kM��sȄ�6���^�A�"gOl�_���L�8VޚB4��c~)�AY�F����D+��zQ$s�������j_�Dnu������%LZK�{(�I`����.K�$w�L3,��RNQ�����d�X�Փ�P���L��\�<��m7�D��Ri�hjϮܺ*�4��OcY$W���mA��4�*�6[Bli��ӹ�s�Am�
�V	��{��p��� �t��H�(͚���ڏ�1Y��0OTNyz����%H��J
(�5��N�������5��'�K7C.����Am��\o73/�+��i�_�6([�����5l�h-}���#��2�eDu��m����=+��4]V�n���n��-�y�ė�
�wR)]�8"U��/BP�j�3��! �D04p��Z/\�O�[i��0r���K�2SMUV?Z]�#��܇��� ��&�	��{�ul�Х��s��ds�U%X|ʶY��z�E�&��1�R �2 ��Ta�H��*�63���k%���s��_������wS����FM��*��	�Na�^���X ����ӏ��q�PH���6�3��������m�`��Hq�p�c|a���e�E�	.",���lߏ��Er�A��ݖ����X��i��}�:��'h꫎�
I�=G2��
	,MΒ�PQ46�QP��n+Nefi��3ٕ	�n
l���<��l��A��a�4>_���O��A^�DL4u`���H���&c���"���|����s/7J�3�����g��l1vC�:j.����-Y"ɢg��B
߬�(h�Ռ��ޞKH⤲Jjw��ڡ.=����К6X��v���(B�G$�q+��!MX��I:2O"�]��@Ze'��L;��0b�d�OΧ���.���I_�(�O�>dY[��y>E=�(��i��0���iRz,G�}��,O�����qbM�h=1�H#0��/��^�,rL ��@8 -��wx_/S�,�#i���"W�A��%�Ɲ����U�<��b� �x��GU�e��]E41�q_l"QV�l���R
t��P�����ޣ6A�TY	�Yb 7�i}���L �%�}���bMYm1Mw�(B����j�Lb��4�������%��ٝx��'��=�����撝�x̧m	}:?<R|�[h����e��>����
$����4���6y�^QC-�߀�l�t����@�p=��kb�gG2t���Tby���I�0�j�V�0�>�f%Wh���թ�6��z��t���4�
ۍ�q�a�@.k��@U�v��l$��T�r��
��X��I�y�R\}jO�j��z��������M���[�r��!p��|ҷ�9���ñ4�i�,��/^3�,N��qG	���KW���<���ѣ��:W2o���/�86X*�H�|����qv�*����>^��)��mVjʄ	�V�9��P�3�[.��w���!_�����	G����'��`�L��,�GV��*�տ���N��� Ά�z�4-X=�k�!�ao\d��Z��,�w����b)T�
��n0���PG����ƺ�� ��71M䳀���V5���>�ڨ"l�Ճ=$ϨÈ�H"_��K��m5`!b��%_؁�L�un�EK#*e�*�u��Y�|�x�y���_�=�+).�Tâ*P�YRR����q�Z����֝w��-��FS�$���"	(��1ҡ��"w(���@WYKB��l����bFY�	�g��S�h4��K������^Z?!o�0<W���x�U>��������lk�A���x���|�$nMM5�>9!�Ƥ<nS
�eK�a�>���2NǠ�����Z��8��h鰡�2��Uf��G�)Ul����*��P�߁�<���3K4�갢2�.x��2�+.^	\��swϩ@l&l����'U@��NY&�b�,	� �\y�����m�'�GE2��f�;��k��v{[�ȟ�]�Xa,vW�VK�����ٞ��=�=��%ͤ�%w=��kY�z�&�t��dv��c%��[�\�qL��\�y�ȁ�7}`����0*��O��
��J��`�^��N$�+��U�6�M,����f��?�mh1�5v�iUlɷG��T�ֆ��b=��44��w�d �em:��u1=	���a<��'8'țd��)�����f����,d�5���t�J���ڵU�@�>���ݵ�5=�BH�m6kUK���o�2K��,��Ɖ�g���w�VcK!ݠ�� *��{�I<�%ְ�ӆ��|f�cY9�_>�&���h�HO;IR$��
dS���	ږP-��܇nnEVќ�-������W�����#j�>U�g�'C�N���_�80��5k������H6�W\�E/H�f���-~6mP��_qf�j�����cia+UY�#MQGT������[��҄�CJPm�lz���M_�|�=�굤��`<fel�6�2.ݥ��u���{,��^}�y�����Hon)�;zAOysbf�&��`R�#� 7��Ȭ��h4ඊTa���8�a��D�ǭH��(6�*D�9�M۝n����
��ٓ�4�ٚ�]���8YcƲ���o���1b��p:�Ж�F>�Ц�캷�l09��M�6.tS7^�K2�J[tEgѽ7C�t@������w7ӍԪY)J��-m����[8(�>�-�q���T�Pp����V�.L^=�=���9��]�j����_{�&���;�����ZA�r�'��7Sc�	� ��mb�w�� �L�T||K�j��f�|I��'^
��dnUת�;�ՠ>�bh��*��)4�B�m��,i����u����րMW��`�Q	eWm_�ݞ�=�ֹElE��=�!ܘ�/�~����10�#>M<�8I-g���/�P�O��a�|��[�E�	,F�]-�=P*�6���s�v�C�e������[P2��NK��|s1NB.=4�	��޵L^�YiX`���Qv�#*h����^p�k1����Y������3��6@�_�Ȳ�>n�q��h{�ޗBW�*Q��?v���I��[��V��v�ATb�d8f�%�Ai��L�6�r�;t�{NM��'�4�1�!��Ӈv"K��ek�Ѷ%'b��
�����4�v��Xߡ�BGҷ;%���K�����^�������e�8*]4կ�0ǶR�"i���˿��4r�}��>�X0�X�p��"jhAL���y��``�a,X� 1�a�o$_{�3: }ʯ�D尌?Ib}ov�	�"���,cǢ��
��o�/me4�+<��'rI}D��
.�n\0���mV�`1x���p�cmO�9��qC��-���S�v��
g,Ii���؉Z9� ]���
d?�n%��$��4im�Jt��ol��A�������;\��z���aw�]H�wU��h�L���"o��l���7�/=�񳶥5e�A	�1���99����|G:*0Cw�FK�ڙ4J����z�:���] e]V����{�w�_��Z�j��h٦		4g�V1�>���K�r��Go��7�#4dX�	__��̓8� �&3z�û�{��q)�i(�a+�Oٜn��w�M=Da�x&��z�j�yk/hR"�3�;J�c/]Uv�xǳs���F&�|VF��l	��[�����rw(��GY�Ri�m��9�oeu�#��`5�h�Z�#}�A2�����N�=��Kn���e����,dK<����a[�<N�@&�i�*�n���IV�������8�6� ��K�f(j���P!�IE,��t]��2eA����1����^���C���V��_��Z��|[��]WqY�j�s4�:�.�2�Ў�q�P�c�N(*E��cR�4K��u�T��#����<́�K�̜��6p�y�����a
�Tu�"��`	�H�=�٦��/���p��-�e�c�c��c��F��m>R�V�`�d ��8�*�I�Q+g«)������&���\��K��A �PG�
 9t�&�~�}FB�,�f	����޿p38�
��e"��wCM���>մ5�BG��V�/\,AO���U۷rf:j��b�VMV	�,-YP��*�.Ai�%R�Gb������u<$�ϖ��j�����Dݓ��Np�Oh�9��k����v�`��8�����">��¡����j��\�JW!���{4>��D��׼���#��IOQQ9&��R#!�@y�D+��!}μ��!˕�jV1@A(tI�-��u�ZA�r�i�'�����Gw�E���ԙS��Q�#�B�9`��%���Q�%D�*�U�r[���!fC*Ah�U���;�摳F3�F��(r�<&�B����F��նC�nN�u�� YN�i"9ܔ�|��i�Nɹ,/כ����R�\p��ds���Z"M^E{�s(��?��S�YmT��^[i�;��劝�SWx��
緼������^q��_0�g[�W2��ZA�8��6�C�Wxݛ}�pk���܌���(�y�l���Zup�{ޭ��1�qGFUtR��SXN��i�E̸[��� �pM���Y9�&�Rxr�����Խ������v�ε�I��x�v~��
������0���߿
�ԶȜYy1"a���k��i@u���i�&�t=%G��y�o��Ⱥ�3C��+�.bD�����%�@t��;��GD�s� ��I-�QWn5R���fw%	����-�`b`��#n-gjю�`>�^U5�k43#���
��*Dy_�y����K�>c�;���a�q8�˃<�/$V�D~�YoX��HH{���� � ���!A�u���"˛�s��61ݟ�ۥw��2���x[�D)V�=�f14��8ۛ�)��=p��7���x���GP{^������/ֵ�o}���@E������4Ms��JU�hk~��:�Τ��ⶌ�m[4)cӧZ^��ｷ�%a�9����1ҏ��B�n��Y� _����,�{x֌��h��Pl�'m�>ZZ�Ct.�U�9l!Vd\�\++{/�ǫ���yIO!]�Q����{���F��쓙&מ���#�[��ӹo����:����g �Jn4O�I�>�����n̬�~�!���C���[�eK��wH�`&��¼rPJ�s�d�{lL�A��>�@.&>K�\�fC�]��D��V��y)����\[{l��48�>���$q�����-u��B�B�~=�4g�#�t�X�1�kE	��z_#8(2�K��f5B����Hݎ~j�L��0���/}Px~�~x��kn���Y�=���f4���x�Bpq]��z�w��� b���ȗ��6C�6��0xc��R�4���w��E�YeyL�̼}8;n%sg�=�F��+qה��w��L��I
��z�6�cu�Oe&��&9�3-����T�\�X�=+[�� �Y睻k�M���nf|�G%9�*��C�b��`��#�������yb�1Rc���Wt�=`˹���8:j�u[�x� �=���B�p���DD'�������D��_�Ԣm$n�wM�4E�qh�v�3�&6�>��_B�ʏ���s[��*2O����M��h�V�˖����n�H�(
$�~`c��j���&P0�������#?�+�
WVٙ��׃�x�V~n�t��0�! P�`�MH\�U���ʞ(������X?�M��o#��Z�%3ғ�j�[�-�BC���ϧ�Ɣ�+J94w��biGRT_,��_����Q2�a�6��0��G�ܟ.���TO�?�N�8�*"7����*�ѝ&G��#�r˴l�%��j	����"��/��c�'_.�T�J1
����g���3e���*^#�k�̋���F�fV�D��$��皩L$��!Ă*��z0�1(��w�Ϥd�)S8Q�Bۓ)@�=*ڊJ4�Z�_���C�����~�d{��BFG�'���qܑ���u=H�
���-�O
Qi��0��[�R��J�
��!��k������#�Ɗ�`�#?��.9`��n�_�^�0�)b��c`D^�M��6�Y����(��vF�r��Ƭ�����>���]���3{�c]봰8E�JP~�)�eX���1�7䌲�e�%p*����y$�q>�Ŋ�����>�dp~�*�]KNಞ$s�=ł[��:�!UL�_{�@����	S��Ė�ʞ3�T�L%rj,��������U�+�T9̚[��f���x����\'��_�~
�-�ރ[��wO��(�Z���ѷ$�����\u+�ȋ3���^�z&%�`�;�pY���d���o�ͭR�@uP�b�͔_�N(�<6����^�K�(4��.����e�Y���K�;]�	C�뮥�]�c@��Wu
<@xǤ�8�ک�:�6\�p�Y�3�z��t�\L�0իfG
��d�{��UWA^&�9�6�'|m�r�,�@�|� �-�C~�]i��5�W����tѹ�.o3-h�̖j>�p�?�1KiB�v������صi-�y��ΰ��u]��oH�D�|Y���(�i��0i�U07�ݥO.o��
�F�}S��-�ɚ�kX����Mo�`��y$]p(�N6=�;gr�8U$�op?xe19�̂m�Yö���Xd�S���6Af�o��C�o��xXR�ꑍ��!רMD�Xz��E���-�Ӛ��w0�ICJ���KS�_�4g�0���|N22�����8�G���h�2�&�S �r�'�Xs�3�%���l*�ER���_���ޤ Ǘ�?�ӣ�����R�������J�����B�L֮���@�W�+����޹��_7�JZVV��IaZ�$���.S��^�l��觾CEB?qq��b��F���Rnk6;��H��s�N��}\�]п�s�+��i�h_v�;�����5<�£�H�M����k��7��v6s(?����uƽ�[<���;����	�
g�S�FǓ���ȕ6!d�z�U|b	K�@�6zZ͔��_Zx����ۖ�<�)������;h͟զ��_�������9�6Fu�*PT8�Y͡�o��i ��	Sb�;c?' 5_GlXo�$j�P�,+^�q0�+Qf�֒>��T�5X���QN�o)&@�M�~7�M�δ,N��<�c�w�l̴"4��@��&͍b��`΋�B�� ��e�_�*���ϥv����E{�ݬ�k����y|�#v&��Ҩ^PÆ��K��W?�\X��0�݂c��t��+��`�����U5�O�-�Ȳ���S��ڙ�?�%�r�+T-O��L����GM?��ՠ�.9q�4��\0AN�:�sX''�����W�+{>TGa�;����;�t��}=$Ce��0,�E��� �+W����Y���kh�*]�WA!�^�����
�b�U,�4���Wўd���@��|mT2�r%!f�\�F�c9M0��ø��ʺ�?@��|�cR�ĥ��uI���~�����ePP�~��1b�fk�� ���-���cɐb�����rf�����8ߢ��&6����Y,��ʞ��^Ʒg���%F�t�=��1�$�+� 'Ŧ�(�<���aE_L��$�А��>T��{�Q���"~���И�y���v�+!,>��!#)�~�_��}{Ӽ!��ڑs���k��!��4Y�]�њ���7հ[�#t�|8���<��"<���@���s�8>>�w�Q�A��)�+Di���P:Ӹ���K�j+���:�>���^8�B�kZD���6�Q?�C���tb��|�K�H0�.jK�n��vRa���iW��B����*.jL��1�)ckv3��������@�&�L�PC�(���V���F�4�s�K7������r|2���s�`߯���S�Ƌu�M-�&�6���P�M�n+�As�1�d��\E��Q�2	C4b�X���Y�FD��[g�*���MHn�w,������dB3�{����95qA31*2S����%N0�����Q�E���Ʒ�_{��a��+���W�q�é��@Qg7�o��N+瓍a:�ޔ�a���h[�s���J?� e|k�l�E'����nG����6��ކ��Ш�4㾾�#樸�Ԭ��	�:h��C*X�.n��Z���i����^�ꨉB68��*�٧�g�����:Y���a�`c���v�c�����eE�ʸL|��ƭ��O#�%��WFx��T6�+���T*����<ܪ�XMc�Ri�ա�W�v2���&"R�/��D�W~#�i��'$c;ٗ��5#��iz�o�:3-��/�PV�uOH������|i9�02��-�m���;*���cX.�(nɎ���������9�l�x�TOLAK$yT��bߡ=�	q�1߼�O-�3���4�n8I��s�˺( ��G����dZ���<ktTN�Q��
�U��m��PC,z�<7@��D��pŦu�Ԇ����N�d�����K`qU%8LTH�j�幝��Nt�~���o	ձ�Tl� ��%C�<g������]�{b:� �}���ɂ����'�Cp�?
PW�\%ó"���{�"�VF�*�(�l�N2}�SȤN�{. ⪠�&��]dR0!�d7#L�*�GZ�֗�3̓f�B�hK��u��KhP6��Q���U���/<{܌�2����`�_��90M�bxЯo�o![�aO����6�9��R��D<1H_Tk>e!���.<�e1���Cr�$bG�G��4�7X���AW6�P��f8iq��S���6N\�X���}g|��E�2��'��N6�_8����kGNp�W=���		�2��.
���>>-<�蹿�)�L�R�>�B�!ÐGn�Zt/̳��d�)%�?�4jJnl���zKm����	6�=|X	�q��@�S��#m�޹� �J��B���Τ�9X�r�'��N�sx�&��c���u[س���L����ă t2$�R��+0���6kvf1�i84����|"�&��������l��J&�B������ޕ���}Jp>�1��e�1�����p�D�������6����� =Fו�tҒm�"�Vc8�Ѥq��k�F}�ް�H��Q�J��[!�Mw4�>4�<sx��٣}�F���x@�wa��8l�Ֆ��h��==����PjW�$p�F�L�P���z9���x]�{u���eEސp��]jq2�tN1���>-Ӆz��D'h��$��ݴ\c�5�#�fT�x�yp����&ީ7�O��\#��;��Eg�]Hi�֐��W���y�Md���\:�̪���Y�r�zDEEch�����:�e��x�pv	Ҕ���MU��ί����p��:'����'_+cJ�ĂY��Mu6N��Pk��)���*Dw�t�z�����q��������I�5�bU��׮�s0��#厤���Р�5<V��9@��_�?3k�
p�SX��+�ٸ_m]UՐ�@x�{����F`@�g�<^'|
]�v|S�lU�gƳ����px�J-�a��>�G�ᩈ�	Ѭ�
3KX��m�:�Zv�m��,�۾Dr�B����L�֓�� B�=�@��M�����'S�7�HL�L[A����R[/h�7w����P��ƓܛV���
�*��s{[�����9{ʳ�7�^��fƪdTm��*���G���1��,���OVx)��yF�\�Op�����2WÈl��͢ZC0{�$�~# =��aL�h_ 04�G�Ox����؈�z����]�*��ѵ>�0����#� CD\��i}˞�v���Ľz��3rqԛ��HDۍ�X�SB��+�"�8����j���8�~���,��#𡦏䎙����yU���Ç��Ě���+o$xU@��϶���>�|)����P�3���|/	x�dX�cb�Œ�z�C�+&��Ca�ܓ�c�{	���bx�ȱH�Y�{'�4��(�״�Z�*�8,�rSn?�T��8��R��C�L���f�)�q`I����d=|����gyƳ�겷��O؏�­)��{(�b��_�`q�g��ۋt8����������K}/;}�ܞ�xuˬ�#�1|��1�D�]�ir��9�C#d9�Ň�Ԩ$�g(�Fs��h��L$ @p��a��	`QZ:�Q�)����Z��Z~~�M4Lf��J·��m�T�Ͼ�v㳀�I7��ø�k��#�M�"l���/4�p�N2g����f�n B�/��!�X��۪�45}՝����h70�����pxQLg�)�*\h���ñ��&Z��7�$*�����#)��~Z�B&�S�2M�
X\7T'>�7����e�H�S)�KT��R;E@D�9����^���N-:u<�Ō	jWq�^E>@��n�AcL�P>�hU4�k`!rMh��X�%��ykID@8�u:N�6ν$pYs���Q6 p-�x0$�xd��d����?�x��-�F�ȊP-��9�<���p��X�v ��7SB�>.��G8�Mw�O`9n�;�u�r�*?.	�1O������X%1�w���������ɾ8��]!@T��b�z\UO	y�&�)X}�K�r9�ƀ<�*	;�;���|ф{P�9g��?����b��&���j6����طƄpU���\D�=Bg�£U�u7�W�
��'�%�Ϙ�iш���*�s�p=t��f���bX�!��J���EV�����}i�i뺱�\!�,���F�7���j��q�{�OSD/+�Y��L[�D�z�/���]�0e+�-;4�/qoO�ɕ�(4�}��ϣ7�L�o�J�֘�od\"�A�S��r&�%�����b�Z3q������F!lp�D ����:�/��Y��V���(G$h�¥*Z���~4^��vB]��p1Sw�c���9��*��:�ֹ�����2@s����.v��b'o
��¼8h��}����qSw�(N�[�g������� k�5�Q�����M��s�p����Ut�:W��%c����'�k��_�Y2:�L��*�M���nGѶ�ؤ�G��u���� (n���g��`��{N~�qY!�Ī��ȴ4*?�w���n����_4�c�����_��ۘ:�%����¶�3�=�+�<]���[�>��66}����d�IYnZ�F'�rA�H1����P�-8ѵo#��.��6�C� ����^�Q��V�o�@D���Ljz��P���S�4���a����	�kA\�Ӥ֚�7���^�Y����q*��n��6�U�4��)H)��qM�H%ᣍ���!/�(X���Հ�4�1�^c�]������so
u񷙇����{�
K��?!^�m�ѳ}��������/�T����Ua�^�|`@�#E_A�iJ>[f!��b�2�Y��;�0eS(��J9q���ɨ�).��o+:�2�k�$X�����ۣ��$�n2�&ڃ�t��ʑ��9�F�����H@
�k� ���4���������?��OgN����x�Z,d]�(:/��w/���B�.-�:�ay��� ����/щ>���K��2TW�Z`���*���yj��,�Mf�ɚ�x��RZ�s�3���h���=�Ji�O-}U�QZ��{)��d������L�,?����hG؝>j�j��帞e?�"߫�^?j�8h:���Mц���_p0f�4�|����'�6%��S~bY�@M�%����aC��ُî΢�ZU�X�Y
�	���s�<��(0���L��˧6���$��Vý���S�3���oABt�Z�������AF�Ilta�Yʀ�P�h��a�L��y������Gj��]�yᆉx��o�Y�MW�a:!����y���]<��$^v���0[·����.�G�u��c��W]/�4C�{�L�r[�FN�f�xȊ$@�i��IQ�2r���4�M������s�_�0 &�t|뭫9�����?�X���u�� �f�����SQY,�m��݂�=�,�x5\o*='-oM�M��ۨ�l	'��@�+*	�N�v�B��Oi�"��n�=�n�j���r�|��.!�k�0���!�ȷ���6�ln�s<@|�R/T�����c����Y��Av�;4a��'��P��F�&A�6��c�-���=,"Vu|��ϗU����@t=�	��u��Q��y�0k�4�	��s��0��'��Շgֈֈ3sy�r�Ujm$�'��(LB�,��JLݞˁ���
>&��̽�(
�{� .u[��ݏ�p-�IĐ}��V�������F�5T����Ρ�$��3Ӂ*\_`J	O@�oxAK?�i[��oo䢨��>g��
{�q��!�`��t-��z/������v���s�0%H�S����vZ�ξ��ڍKBy*��+�n/?bT�(/)�;���P�j���I�h�WHT�԰�9�[Z�:)�^eu�L[�����b��b�����+��cH|:���$L��Z��O��d��3�Gx��gQ3ݢU�i�u��3jk^\�1�� k<�r�E7]~�t��ÚK���b}d�>����&xx�Z-Tk���ZacI��ŉ�X��tա�1�d<��ָ�t�qJ"_��3�����8��������3gtNwk4��}�������	��4��iK+�h���������z@3U�B�B�������	���XL�fCzj�ޓ<±���Nf��#��%Ƞ*dp�)�V�+3�w�sy ��б���ۡ�}�J5��V��!�a#�<�"��vv��Z� H���H�,�Dk���N�0	B�}X��n�ݞ9�yK���^9	�OBM�H��]p�0��� �Iм�Q�$��¸��w�XE�@��-�2l����+6���+H	1gg+��q)@��o�K��㉒����� �*���	�w��/mgڹ/1>FA�ڃ�o���~O��+�NL� �;�}L�Ƴ���50�l7��&��h".����߿�Um�ˏ��`�(f��)���;Zs�,x�w6枎�3�j��ZaWN� ���dsGP��`�`���t#R<勉�5�<�!�-�����B��l*i��6XFZ�.@�$�+�QD ��~Ѷ=��x����}|x�����bp@2И�$>��9�nDܒ��%&��}�j���u��}#+,B��_��J`>����G�;Q�I�殻���w��az���i(�B_�*`�>�%�6x��W�$�<ʸ]��Jda9#�� )�`�
����D;�n��\����*I��Y.G�����4� ڕ�¹�b��<4���V��@�����"�QF� �q��k��g��M�=�i���q�"��%f �9��b,(� ��YG������2��c	���fr��	�k�B����M�K�<-����Vީ���)�����mߙ��9�K�L/P[m�M��J����}�M*�s�~���������z�2l�ڤf) >�b29��U�Zʳ�u=dġ�#/V_[��>�p�*NsS��hi.�����$qn�*����3�3��'Q��}v�s_�{�	�~�|��x�SV�G�[��(6�(H�������ow��ssv�L�斤W� �l�|��K�FO^�n���h�>��o��4;���s��`J�}9-��pb:?NZ��A�t�x�3��~�r`��s��jF�!vP懲32�n�F�5��$9��)X�k�C�,E�|�ƭ����E��~�}�:�p��]�{�z�in���$�W�a"̚���ڳ��axɁ_��²d�p��$��k�K���8�pw�Ε�&c�e��&����V���-�o�#��P��9�'`�%����y둁�P�F��@�u�s��$��e��j���x�����7�=��� ����3ȟ&��uX��s!-��9I|�
i�ɣ���� v�����4�+��n5/g�mX��������r����45��T�SH'��h1���9�`{'cW	�e!KL��Ǚ�Dp�$�zZ�_ �`�#%��;t�͛!�j�S��V�nN�������}�-�#�gVDS��߷�b7)PE����Q{�2��q7�ڲb���t�ͭJWTۇQ����9���t��4� ��<�$���QG�a^s[�Pw��A�i{���<��&��	�LvfTE{���x8W�C��;cŘ���6e�Rf��$����9�)����p��H�:/n6�aWR��)/ŵP���M��	˟�HB�� �&�-o�{o�	����~��^��r�~���F��r>�C��y3��|�w+�ίLF> K�ڬ-"s��WQ��G�N�
i�K i�-�ʉ��xb,�#~�qt��'��'�_��ʜ�2�O@��?���lz����ϴw�{����?X���F��7ٖ���
]�F��\M����y����ݶ�����F��$^�8����X6�_�?PR
	F��h�C��Y��h�2 �h=@=�D����?��� ;�*yZr�MQd{6�Uj��� y`1����&�:�����&C����+u�X�����Jd��6X�e��li����^	����E����wQ-�13h���Ǩ�n����%J�nݛ �IYj��U�4O٢��i+5)g��]	&�����S��5�_]鐳m3����x+�g�]be�9'�I*�w8,~���m�w�mk"z�3=j��1������8� �*�|�IU�>+K��qZ+N���
n���K��%�Q��k9\i�V6d���p��j�Lc����Qm�4D;�=a@��D�.���'���$Z��ң�������o�\LR��,��eLFg���`ڜ���-p��[Ǫ���
�_�M+�3�\d���D��M-t�������S���O�d����oٗ��W�9��oN���<@�D�o�R<,$?�e=6�~2Rd�]!�A6ϩl�Ȣ-*�����r��+/$�wf�f�E�霻N��|m���f�"i^�`�ц{�<'�
3��ĳ����`:T��0\�F�$b��וּ�ktzh����u%��@��ᝆ���WT�E�+`p�BU]�4m��śD�y'E��'S��G߭0H67Wy����A4'V4��z�n�x�c�a�R���O�3���C,��V"}�yv�_@����G5b���ށ�_%�u�1�T�G�>恺)�
����߼�+��4�b�Zr~����)��C�1�oMqA`��PE]W�{NNn�� ��#;+��!���q���J�~R�8L�)eFH���M��pn�0���_jt%�ܰ/4�=�	��	���#�\��J_G��H��l	 �H��,�:D��9�܆��M������@(R��9�n�H��Cm�3��{/��"�U��i`��}�7`,e������r�ԯ�c��#$�����ngz(������y�I@گR��w������
��]�i�Yۛ�Wmʓ���[y:iØ�����X�H(�g6��\[d������,�agVY'{4����ws�f%�"lb!�,L����E~}rc#�72h;������vঁ���w�;��!k�o,�>a�ӹ�~]@DɧX�Gy�*j5�8���D% Fx�UR�4D�%(Y�-���{?�v��y���<�1��c�)tΏ��f�}�sp]�o+2:a�7�]����a�l���O��������I��\���3��+� ���C� κ�4Xmy��i���˾��j�%�2L�¹�+�$����*
*+*v[I�Nn]�P�F��u��r!�$6Ѡ����P "��zS�S^��C�U�Ɍ|�3���,��,x����!�z�X��i)���	�d�c���E3G���<�A�Z!SJ�!W(�q���6Fm/
��+)��u���l��b{?Y�W� �!Nl�_6q�1x}�Q"�S6,���<�e����\]_YC7�g�=��Y��������3�<[}ne�ʘ����g��{>�j��J!�+��K�:��6]K��@�I�\<��|'S�Y����-�[�#	�_`���Y�W2�O_�?��i���Iu2��,&�v�rn��'��d?7Ig>��|9�eDo����3�H�����MD�W ��2@�"0�z����c��A�\o���z�CN��f]��VA��q�phʵ:01n���bdE4�����~/�9H�x��5ՔW���h���ì�������@C �%�T����;K�YH�B���]����Қ��PE�6u�N`dn��+
��-�e�V�j蛹�<:,�Dp	Vd��� &�����a������[�H0n��wea��`(9X�!H�)#�9�Ԉ[ ���Z��om]�����<�y�%�֯|�����s~�|F./5(#�[+��������������9܆��Zۀo�e,�oȭ���C���E,X��BD*wa6���Z?�ent+�  1&z���,mZ�&�"��|4e��c�5�'�u~wn�v���������(�G��1I�	����
Ye����i"�C�P�8���J����l���&��+���΂AT?ٰ~[m <�Xk4��U���jI2쿋j���Ph"O�|�q����+�KT�ne��iif2� �&�������<Q]�o/�	΄���t�����.JF�����682��D|�ZD�LX(G���#�;=��ioza �J͒;�D4���A�2 �S�nE3��F,��ץ�9�lo���@���쑩��>Ep���Uo���i�_!�3#v�]�rhc��O$҈݊¡2lӨYBׁ�qA�F;��v����G�(�K�3ͩ���S��I�L_�^��(�@��s�ٲ���J��v-��J�_k�'�ǔͿT��V��2�}��y�6��`������Fcy���2_?=�2�_
��C�|��w���c�Ϟ���ƻ4\VQ���!��:4�:dق�� �U��iB`B���٨dPb�U����q���:��o���!�@�i?q?���~�O0���CJ$�D����hc&��&�Y���p{��K1�����c��b���%K�A&⚙=k#j��M9�����ݣ���5Y�h�����2���g�e���3ǴW]��~+��W߅i1q�=�o�m�k޹��c���6��	f���ޭ͈v����=i
����f��Ã`��W�-�l�)�L��A�Y��[��O�1sT���4Ȋ���Nf���k��Hl��FP�!ݬŉ��n��1UV'�TG����϶H.wiGI�c�v]]YG�����(�-'�ށ�oN�%5<vQ`�)it�^���tzT�iN��t���6m������>�\g!G�ǣ�X�惖I W��jp�������ę	��	d0'z�'%��W���ӘC'����A���8�Z���#���%?��j
��Q�?�ܷ�_4Ӂ�V��.���ƾ��੬�z�S�d�\�yHȨ��%̃r��+�
���VUUf<�!�*��J�%4���6]	���偻����+�Q�j�sR\�Id��9��oh� S"��]F%��^v�ls���#��B�%���=��qj͐�
$�`��;z�Z�?C���R�U�YJ|\^D�%|���:-��MV�{����x��P^��d ƒ7oB��4���Yc�W�����<4�,z	լ̴��b�m�}^�?�ͅva�Q�I�~��ON5��%Rbz���5�ų:������A�m�Do��5��MkKj®�&rȎ����6t�v�h�ֶ�k�ːw[Yg6�q�&ƽJឆ+GG��ύ����6���N3�[gI��隨���@���M��T�q���i�}+W��HW^i�x=�'�ފ}͸���+I�s�C����9��� �Z�_ ȼ�	"�vvdXr	GY�H8�����Y�<2�h��Vw��2Q���  �@�|^�&��f�w���<[�	���q?L�o �@�[��.
���)=j`/d
��d���N�/Q��7�8a���1���'PIc�mQ˥�\h�"�/9�at�V}�ؾe�� nv���BǼ��HQf0әs%@²?Af��N�� LC�0����l��j*�	����on�0k���E'\�+��>9����9O7���}�['N� �*d��d�wp�1�U�v��u^�����?��G:�7��d>'��~S�B*�B���-&+�7�7Z�'+�[Y@sٮ��c����~������֩��n
7����9�NA	�֨j�u�/�{t'�f��"��e� �N�=�1���s��&
v5��j�:�yv��i���6}҅SѴ���tȊ�x0��0{I�1~�����I�÷���V<n�.��ge�����+�%/����h� ڷ_|)2UW����4�k:�S0�Ԍ���3��'t����*�i7C:ޯ�b"��e#�fͼWy�9�z���	<�JC�6Ï�\�2�F۔[c���6��mk��<e�U"��n� �O/��<�JME�5��"��J�?0L�����
������y�{���hv*u������X�g)�����cFf�۟�V1#�i��abyA����މ��������K�Ԉ]��ϋi-1����pٚ���0�®!��O�<�����i�J:��R":OW4�A�!jPb"����$&�)�E�kF��b�{8��JԒ*E
㍫�Ƶe�2\F�H�S��ښ�����d�m��=YI�F��Fj�iN)�:�k�e��V�訢�e�xn�4.�QQ໗'��g��;Tm]�m���,"����w��L��m����Rs�&f��^t4���+j�b�k�U4�է���?��I?����/6�G�v^<^��p!4��rL���G�O�<?���u�>i��������b���*���rb� z>�'6����o�X�@�i���h�_6��+�L˭�<���:�.54�RJ,0���3z<\������;����p>l�����~�CO�V���?��d"�c�v��'����$@{�2�y:��zߤ�@�hu�V���i�0�G��qa�˂�weϵ3���ݎ<q����6�w�Pq��W>�S&]5��p)Q��+�T]��Wޮ���zƠ�ނ�����g_��I�����ߥ|f[�l�t<�.~��չ�Q[b����9�9��;dy�W�-ruWs;{��0i
��@�K�g�Ij�3R�ܸۼ0t8#r���hw�S3�~ �F>sh/���ǤM��)�3�sy�!nʉ���V��6d|e�Y�e�\����p�oh��!�ϝTq�����+֮��+�/�cuL�a�9�J�ݯ��P3_5�2h�
Z�"SQ��ґ/�X�<�����U��2�Պ��,����5��c�e�̒
�*������F��m��]F�*�Ϳ(J�k�� c��p�H�-`��b$%��ǜ�(��~�����Yq�'�I9DS�ź׼�ٷ�.�`�^>��� k���9;��V<< \�ĭ5�J���:*
���;��Ak-�1�۷�a��,�����?���^��AŬK:�\0S�}�8��4@��/�/����~��Fnޛ�h�E|W�C�A{h^j�+�5��h�)�&	�ߜ���q�C�2�U<�CoH�+�[���ɻ^+HXq]`A�[��< \�����]��<��W�9����y��j�<q	Dg|B>v$%�+���A;}�p���VB'%E����.cflR��9C$`BOBsH甄`��a�I��
�A�A$�V�lk7�W�)x)�����Z��m4�}�r�("m����9!܀#k!��'��`�#4��.�D\�]Q���ӈH`v�e�FeW�A���o�>P�G�u\�k�
��������H�Kq�PS�}L�Ng*�vU�y`�5K��(�al]掚*���ࠁ̤��q6�$T8l�h��J?@N�8��ZG)���Xz4V�v�Nr&$���b�����n����`���~�`mM���^Kܣk���j�z�Q69�p Q�IB�p�&�Gřv��|�a,�W �SY�!)�	�k�@M���1z�FMm�D���;��n��C��QܝR�6�_i�b�SZ��x��F4��6�~ZN�\!��f�4U�4wF/�E�9@{�_ː� Br�=�諭w����]��ħl�Jb��DB��^٢^�>�3�����y�F�� E�o=�؅'*Ֆ^n�k�t��Jr�ީ��"���E��z��4��J
�#��E�	jn���܉����)LE�z���t4)y�h�9P�$��hG� q�ܴ�Ѣ�l� T��!��sx�"�#�5]!��`_uAS^�M��~��bZ�4
K���T}I���YQ�n�s=�L;g� ���x�q�h�T�b!Lf+"���_�Yy 6[�3L|c�({)YL�x��� D���X�R���G]j�^O���8	���Y/y�׮p�9*Jpx�'n��4���]��`L$9*�����IiV����,���nu��m�R� s��-�W��#��c�������T��I�4�\7]�'!�1��hn�ƅ�krϪ���X5��>]�B��.Ba���q^��v���O�x}r\�,)��R6��^8h)8_i*�}֞_���8�.���r?+����0��J"��R#�� H,�!*��9���Δ�$Ù+d,�ap�X�q1-ɺ봽�_�>�0�Ar@\�I��le�
#m,���|�E���3������N�[Ċ�f���4���m4t)�bq������A��
�w���������vm�:�I�
:���!�����d�#\y������ �ܧg�2�oP})du���KW�d4m�����񟟦��m�@����J�q��Oч�PV�w�0�?8�ơ3/�z_�,�=�c�Uz ���`SW�vu�B����yJ�tڻ��cM�hL Qչw@k*?�H�����-��:�HK��<��T͸]���*jDK�Uq�(ݒ�]:�ٟ/�&���T�:�}�d����T��b�f[�닲w�6����	�0 X�q ʧ3��o���2�� ��W"Oů��D��(��W��|��� ����<Lq�߈��:�HS*�}'�d)���&��F�@b}�[$�g��#�Do�:�ھTl�-��2 �F� �$i�FK}�jL�L�!�aM�2��N+09�w�|���=��58�J0J]�o@V�N���sI���Zf��yѩ�Sڪc|�����aa�Gg���Q�I�j����2v?-�%*�,$f�g;"ۧ�&���vҁ�"���8�8����3�)��{j�0�Y#���gCܱ&�I	^�w��B�~կ|�C�.�첈�{����<���/q�<+�7$y��bg���l���X��nwm�Z����(2�F>ț���gt+|6&-�h��ɊZ��D)�`jƜq5{u!\�jH�+��
zc*�?,L�����Dmis6Ѕ�=j#��|�Z49�vq!Ur���{ͬ�_����,-g8BdJ1��𐺈k!� &��έ�:��u�'*�6��D?Ob��	m�&j��U��L���`��Uۅv(e��u�Y�"E��O����"��/K�bxb;��;������i��f�8M��3���̰�,?��U��G�E�:H}{�@eu��R@�ƏٸA���c3ַ�~!0���#yW�#��qA�L�B�F� y���R�ɞ� TN�y��zyu�l�Хu-!�ǽ>90��A�����!I���;��TC��Ԡ���}�������Nr���N>lY'f��`����.�`Y��E��m�)�|fe JǷ��XG����V��g�$�3;*�N��:Te@+�y{�VnR?�:P�P���N�U��Z/�[�"*g�Xމ���w8��j�B^�0R �T&d��_A�[��/���R�Bq�%�PW3U������(W}K<X{�P��z^�v����ە�:�_vӵ>(�^yRU��++!#�`gg�^v��o��-��=A����H/��9��dϖH{x.}����~��J�hl��Lim�:�����pP�34�S��p
`���%������Z���ih*���ьW*��qD�����Րƈ�@iD���abW&SD��o�C��&�әD����Y��g{��Յ
Q�J>�a�����%.���!6A!�\�Y�v���3T#�0��	y��J�C摿��-VF9.��b��XC ��Σ ��j���d�cQRTA���T�J_m��4\�Q���Õ.qG�B^T���	�KZ2�0Vkb�}��P?vb.p�{�#{�=3��t.�n.o��%+�Z������%�Pp��㸃Y�<�X`�3+��q���*�3��D
����͠\�S��-���k轾o�M<��	���n��m���l^�p�ĸh�&�:?f�V���1&���3�
�����L��ܿa�`>y!���v�0f�Чw�A�I@�U�G�ǵr�cw�����9�Z�}؃�͛��$B�����^��s���l�d�Ƚ��N�����MB>���V�	67#��j\�{�i|z��ot��T��퉢~`W��U�ߵ���bб��u�ɫ�~�����8���q��F:��kK/���2���d�?(�9�n�ǆ�,h��O�dB�'�JQgtl�B���r��T�bY��;�h�<�{���j#=��
�KMo��7h?�ɔeИNRi��Q�9�>y����F׶� 7����!���p�`/�d�)���|E�"��lAn�@�����|��3h}H�j��;�cZ\CH��D����fM'�pqkB���b�d�bwf���}���μ\z��@��ʚơ�L����Zc���s�M�
�>c�@*>p$�g��J�~w���P��-�QL�IC�y��y���-�Ax`��QN\{��Ľ���Q��ń�<����f ,�����7r&�/�!��F��rG0j%P#ԇ,<���F��^� #G׷�(1�JX��Y�cVE!�:�H�6@o������J2�ͩ��AځDR�����t�7��n��i�"�qv5��g%�[h �M���1_G�+�(��a�/C��ה|�	\�3UKa������z�������&�~݁]� 2QL�7U�GQ�	Gn��1�	�=ߠ�f�[�6��h;��اY��j����d���M?q���"�ƢTL�����涡��Μ�p/�:�T��
�"t���@���(8�P��v���/|���ɀR��Z��s��ˁ�I3�[?Ȏ'�^����]��g.���;*)e��4�zf��w��@�x�#cL���~�v�f;"�i��};��n�� �)������^t�*{_U�d���)w��ЎC�	��խ�w���jMջ(8o��:p )�������H.�h�z�px�4��al AV1�%��i���)em�Բȁ:i�<K�0le(n}����N�"T���m�j�K7`W�?K�{�i���%f�J���N��q,�LC!@�5�T�ʯ�y���NBP�����5a���ƙ�P��%i/L��[�ծ��6��P�߅eo��j҅��&�?��ʻ߀�.l����߈6'W�6!��v:��N�h�)�$���EY�" v��p��z	�T������q�u�L�����|�L�k���U��7�[ڋ	�H��.�o�h�����[�X�9���-B�m��"�%Үy�}(pt��]����Ve�ꆃ ��\�p������h�{=R�%���%�9�95t%�t���{�A�r(����ӕǨU(#;AD�B�RB$�nS����w�s�%D�pޠ�w.-Q◈�a��_Bx~�� GC��+}�N��z[��]� ��|�}!U�Y��MnJJ�56�1���l�J�B�WA7��jZ�D���l�bok�����g'T�h�Y��<	.|����K�@��b�P��ۏ�;��S��8:0E�����-��h��:bDv���>��"$T�����;b���L�<�ɷǉ*R,�Kc���Cbk��DM.���H	�������%e���uXKR������}�_�ۖ��`U���b�>�pBK��*$P�,dY�!�5��U�����j�=�jPA�Q<�.q� �� W�������2WdT�~{%0�U����4����g�`XG��l� ����e���+Z��¸�:�5H�Ő@�ϡ��.��s(1����\�jƞ��:`��rx�!�r
���`���زzi{4����7'�$�5ȃ��n�������^��x�丘�?�M�l���}{W���`u&�4�F��U28�t�s�r�
�!�h}�r���}^l;��;�bE*��_.�T̳_S�pS��C��i�	ܫ}Sw�N�i(P�O�m�����xIYpn���[��b����C����#0\�rB� �`0)X�A��/��s����ڿ�*V~���H�������/���
��a�W�<:x��
*�w�g0~x-�μ߁�$�K��j��ޛ�ۢ$r�9��I�7� V�q��y;8�|�r_�q��ޱ١��C  ����X�����&٨��^�~>��g�Ԟ��Jd~pш�Dҥ��60�>��STΛ2T��P
�d�-:�3'CS�Y�j �G��MYd���3�`��uu�g�w�p�{�o����JS�l�5�4}�iA��g�[���A.��K�p:N([Ë;�9[Q��6p�:�k��z�FMR͐�=��pRѧ"ɬQ;=ی����w���n��j/�+-�n»È�HN�<Y��9Z\
�f���!I�/Z�j���x
�+�Ս L��l\�p����Z��'~�;!�{:�ԓ������͕�D]1*�Ͽ���2)��T��2��ɇ�l�#���e�n�֧�B����[l��?�Zz4���W��@��i�`��A���[1��]�A:x�Tf�aכ���P��xt-�Z�+}�C}&����jRn�]���N�9�puv�:��R�#��m�g2��C?���t}n��L��,���#��h��~�Ѓ��~̬���cty�e��Ԭ3&���׫`�	��suf�x������	J�-�h�r�Q�;x�(:���k�{aMD�48���0M03���������ć����$K�4��S*sj��j�S��x* � M���ï�� �_]��S�ѥ�~\�>\R�4by:֋�I�Is�< ��8�b%ܥ+�k�����K*AA�#�!��|k�NW\TDjSU*�ix����݈E�nAő�$x}č(.Ly�k��vPdj�N�m����>�Ƚ�=���� 򂊟�d06.����e$�E����[{������[�5����ͯRS�Ź��I�1�E�-^��h)�di�m�ֻ�6�OҦ��p�,}�ٻg+0�^#�^�C��g�V��,��&����N����_�6a��o�X\�� �H�����ډ�/���w���9�$ox-Y������/�+5ߛ#�sd��^��w�`Ո�Ņ5Ĵ�a�� �ۼ/Q�*�=A}m4tJ��*�kJW�H�
�Z������ ��x�_��e=�b6U2f�)���ų5L+o�� *�������Sb�n��i�C�4��S�iTWD;Zy��~*Ԋ��>9q��%;�-d%'�OyV��)�ϋM&�Tn�U��~��8�o&�(��������Y��P�C=8�{�{�@��sbO���h��_`
o�˒������z�+nb��?�n]��_�Ұ0��f���mKԅ�SڛX��U��R$"�~i(��@��o���,%k��p�\G���iQC��b~#B�OD�� #��aT�p�c+���:ߢ�z"7��G?�<�f������ލ�ԭ��E�X@�CO��:���٩w��8�BdУ��jM���#m��Dt9fٰG�/.� ��BR��W��d�'=�u�@�oyk��V�g͠�.���£. ����g������g��rqѬ�8�������?Үx"��I/�r?�4z8���h��E3I���fT�x2qE�s���a#����"(ɜ��������Y�w���F��٤J�T�E�Ū��x��>$���q��d� }�����2{����8{��{πK���c~�4����YTk���41?������lZ����P�o�}�?[+��FhO�I����&��z�k�X�*B�Hs��zh�:����^�K=<n@�w� g~�X�.M؛	��!�i�t���E���h:�QM?([/�h�Y ���M?Ԓ/$���&a���3>���lok��hP�J��M�D�1��
2	����4�M������Fy�^��ȅ�E�fɛ��^�'���;�N!<Pg�e���_�#v��r�w���,C�O./EA� ���_�Q^����b���n���&��Ol�w�I��$*��y�n����U6�Z���*����IN~��&��VЗ0ɣ�07�����z����q�Z<ȟ��gaD��Y�OȔ�kn�|����
QS����)S74j�1��B1aZl�#��Eq9��R�S't�M�W)~�5 ����7��}���"k���ϗ��ร�!b����#q�ÊO���<��(�|Sj^��HK�\D��M/Sv c���`�S1�dL��%��C�\��ht��g��ذR^_�%SzeȔ��&��|�d㣕3�z������ENdc��#�3ㅏx�I�Jj�R�%=���je�̈́����"`�x��m�� #�OO���/��5?������W�А�~f`6;�fW�����+��~�Jf潓� ���!(SC%���f���E�ϥ������N�j��VAeH��6�4Θ���2@�X�>�Q9E�ϫ��'�N�~���V�e��*���Ј(�%Zu�s?9��~�I�E�EF�IL�Y�p���IB��CCuf�������S�}{t���7���5����
Ŕ��]�[��Q�z>`´=�ɤX�ٷ��]���_\���O�Q4`U��|��0�[�!�T>X���Z0�����B�� ��:V��Z1��Ѣ!�49�d����[��
�B� Oȑ�%�t�W��ߕkS{p�>K����_��.�ޥ�z�FS�\�]p���KtE�w�ƒf��t���%#�t�r��6h�O��<xN�NW��;PX^�Q�'C��돀�~$�!������R{S�(���JqY<ە�aͅ&��-��4��y�5X��	��\�T	���R;3����;�A�����%�NF#mkAhq��υ�԰���s��*T�(I��91�ds�����\�����i��ɨ��29�'�CZ��T�W�x�Y1�q���rT��Xԣ�l�m��pA�}6���i��:K,�y��LF	�0`��Sd��LC�v�(�mtQozz�$��P�.lǼ�o!�M
Kj�ue��0��dҲ�T\�ߗNtx�Y�[����Q����nÖ?�l̲���|����ƈ�N4c`�')��XŻD�r�w���ԗ��
�ϫ/O��ʍ��׌�<P��^ZR��̉�e����������&Č=@����ϳ�f��
3�|g�����C��<n��_	0�ȱY�9p�Fz-���>�!��a1$?����	:��$%e/�_CC$�;��{7���	]:U+O����'����>��l��uYW�������0���I.��_��%���ű	�:�Fmw?���B\: 1Sd[ds�Pb���Q]�=��А�"�+� �����֣��I7��O�QF��V ?H��C����g�I@<�$���g��L��]"D$���ݝPr����
H�ʏ[��͗�.ˤ��1^f��6��SY, �0H#"M�	Ԭ���zϬ���$��~�𷟝->.~B@i�$C1�����\�&�rn9\���ſ��:N������qH�/�j*)�_��OY�I:�R}\/���t�K︉P��X?%(�_M0��腗U����h��	���.�-��"���ܧqA45�qR'8@��ض}W�!)��!�3�� �u��=��R'W��ڤ�YNRO�sI��2;BwUn��&���~~Q�)�.�U2�-�pL9�#0Y��~�������HU�D�he�;b�3���-v������a$&�>L������#�S&�g� 8���{Q�ϖXLi��VU�e���+9�3Z���Ҵ��|�� �R��L�1����|-�B���2�5PH-n9p<����1nv�ձ�GK#�'�s���}n�KN!�q��Q6�\A��o��\.�������o~3�v�����:�)n��m�K�pYW�9�=M/n���&�C|�,�(M���щ6�[����.����¿S �uĘ��=���4�2���[yr�I��d�!�v�k��2�Q�46�*,�$A�������!xWdFB���)b�LE&p�J���IVe�,gC�L��"'P�n7amy�o�tNܞ���i�	�Д�6�X�QA���o6�2�s��J��¾i�A��\�L�ÀŻWF�`�"����;�	�5Ӱ�,"�P'5~?�����Gr��΃y�m�g	vϸ�q_�鬙��'
�}6���יs?�ז��[�&��:�N�*��]�Z��hZ{!�p�J���P1�\�펱�����p[(O�TD"j[��!O�V�'��B�6�U�p�w�hy̡;1��oڅ�ɭ?�����Wr(�k�{���E�<-�)���:��{}�Ͻ���Oj��a�RkNC��,z�
� {�5ˣ�ɝ���t=�<6)����I����D%�O�7��檡�
d���=�Tc�-Q!�mz�ٹb#��qxjK)�KkkD��\�u��/��@��,�L^l�tER���ǗB�
�he�v5͘�͊a�wf��� �k���������c�*~|��� iR�#6�������8����'[Y��d+�����a�)�N��~ߔپ�����s�A�ϋa.��=����m۸4wcD��z}��j���j8H���SFu�>��lI��F�6ӧk8��V9eN�	�At�`���N�P�<����Z+\b�Qm��J�e�^d%3������R�-��ɮ�R��Ѩ��j�*�c�]O�&3����"U�H��C\yH�>R��r��5G�f���J�B���p����Bѻ	��M�D��j��)���ce��Y
����R��Uּ��ǥ�̦R�$a��T]�<'����P�)°D�*we+[�ݢ؜�F�;g�DZ4���ӵ���O����/�\���N+��N�hR­�
z��B3b.76L��`�; �i#=OJ b��UCN%���<=,���2��t���]qX3�(xoj<��3)9�a��TuS���{��}���\��b�ymRD���2��;�=�L|,�];�0(���l���WB�5�t�b�p@f�����L7@堏��e��X��~=��Ӷ��6��"��O;6��U�H�f��m~���¤�ν�z���Z����O���~5jH���g�U�]�������}`@b֡�sP�"���}WX0�G�n�5�ؒ[ʑ)؞~tZ��f�AJ?C���ܱ%_�D0~�c����31����N�G�v�h���-zʼ}ͺՐ�p��~%�w蔫�7n���ONA�]�{�ޕHē;�vI.n/�.(���!&&�GiD+��ɧ�Bh�ʇ��ʫ��A��F�k����.��֝T����T���C�b:��.�9�f�kl� �d�0c�$����k�^v1�Ⱥ�����d���{yW+�*ڂS��k�a-H2�P�$�A�ZH�wr4 j;�g�e�[b8U|�l&�Dk1�h6�m1��lP��|�ɺ��@H.�����_,��^�\���䠏_�E�:搖w����VJa�=��R#y$&�~�#����`�Kn��R�Yj��J����.����s��G$��I��j��u/ʶ�y,D,���Yf�V^�i��2[���C	���+yҘ��qs�6���G��3%ɐ�C���iF�J~��CX�U$؇׽�$��y��H��g��գR��0-�}ϱ����?���J�N�|��o�̘�̧��l��[�#�}	�"�i#�����8�oP=5��E�
c�잠ԁ��k��<5l�D~�S1�[ˆ
�;3iSS��9��1�q����ر�@��{n���"-rI���A���x^2mżnI�S�GCGh�mb�"~�cy��w���=�L��սE�Y�Ma�� �:��U�^~�g��e��r$�P������^?�%6�D����e|�����K!ʱ_Lx��gU�	}�՛����F$�Ip��nͭ���������m�8]��s���:��������R$oXXj�E��<1bz×=�ϼ]�y<�/ǐ����_� �o:@N_�-��ǉ�k�B�rJx�H� �]'^��f�hi,�gN�����ڈC�ruU�?$��\��m��$<o�D���"�e*gt��Tֱ����b�R4��e+��!��+�z�!#����r�� ou��!�#c��|�1���4��߱��y���aY!�w�tޙ�Z�A��R�I�:m28���e���(�3n�uȝ~��r8��b�顖���ŬS��.���|�d� A���*�b�E�j�$pxX�B�|ȽX ��� b��`�@�8����Q��|��1�2j�j*W ×疙ٱ�+v�O�[�;	W�H��(�E�q���k��2�Mu�L�u˶�ˎ��o�ز���X�/��ޥ7�0{E�?�O�<�4h��r�8�*YXS��w��F�r@�li��2e�;D�k�y���g�
��]K�G���v�i�sN9n�{Zz��5i%�:���"V�ӎp�{tC��"FS�	�(^�mK�ib���Hgn9e�W���Y�
y{�.{�?�w)���46{y�?�ۏ��<[7#F;� �R�f��Bɸ���3�y�C��fIpo]�烰Բ�\%외����T�.︨�����y�7�f
�\J�Q�|����j���������h�K�[y���y����)�R��F�f��3Q���dEl@,��b�|�l;�-�����9"�
̒����K#���)�h5�Ω�+l^�h`\1�ϝ�sn������}h���0���gq�'�t�H��Ħ3Ll�qd[�K'���,]�k^N<��n?��O��������X�O��[���t�"����]u݂�����`�N��;��o�����(�mf���OI^_�7���s~Ԣ+��ʶ𘑄�T3�QI36��\$���cm��8�R�IR�,�έ��ÅH����,����s*��A���ޞOBS&� 9/ڡ%z�C�w�<*�.���5�X�鲱o���A ֞ N�V��	�*�j�h�gAd��(�Xi,n޹��"��V���0��kyqAR�|�P�9�Т��sd�;6�gm ���M_��T�E��k|`'�d�!� b
���|0��[y�C"�C��4��"�c\�:��a��O+�n7���^�E�������-D1�gf}�;�ΨO|����-�{��P��g�U��ypUm�|`*b��;��'�]�r�`�v9�[{£|�BM��B�ehH��X�rˈI;I�1{q�M���r���!�����n���{��x��c>�
�U4�6&b:����	�����7�;�G>l�86�W�U�U��kL�ꘔ��,��!4�h��EԸ��'r���3���^|${�"���`:�n��c�<��d�B8�����]�i"J��;��2ɐ�ɃI��
��<����"N�#�r��2�+�صM�8}�|�����AF�,�{v������6�����O�]/�� 	�'р�{��I��$���7j��tP^���zރ[r����R��/跎��?�zx1��#y�sN��G�	�{��� �Y<����a���nb7Om�9��>@�UĢ��f�>�]ع�����w�(l�2kh��iɂ'�歁^��)���,��a�c��e��]^1 �N�{����E��Sk'��Q/�`&���=�&�ts��^�˦'ꪖk��8�]p� �wJ���#�{�}w�ǰ9$W��.j�ǯ�*v%2�+_�M���:�?�>��*,�!̗���:��)!��b¾}���iЀW�5@�Ȑ� �������CV�TX
x�C�ӛ>;��V�,�c��9~�7E��T�E�OA� ����ϱ��+�`�nSR�zK��$:1Y�� %��2�rM�x�fȅ���,ꓖ8^,�|��n\$�&�&�m�W��&g�L-��T)["n��Io�+O߼�D�_���<���4���7��⥋9_��c];���W���R1j���-�~��]�h�u�X��"�4����y�Q��˖P�#��j��lt�#� �x�ҧԘygv `�g,�����<�6W�ik��X�(��~���i��V!+$�c�.T��WX|I�6�_�Zd��{5#r�rngm��+��6��îh؄|Ȋ}Gy��}q��F�� �j�r�'iq`��UE��BZZ�
�������j����|S[������%�C5c
 ����u�dW���&u+Sp��ь�O�By���1�f��)Z�21"�}�O�ygC�����%�@�Q��[U�ɀS��p��YNb�k����wt�<�~����x�3(}Тl�I�:fBD�c%�ސ�&�|��%T�	]�����i������{#u��XT�1����&C���r�az�J�J๸ ���Ϯy��w��J��U���v{O�V�t�N$r�~�Y�1<>�OƮ(r������=��f��gȱ�T�fx�'�g����{��#"���l�Ң%�����],��	e�9C���Z]�Ӈ����h;�����.\�֖	��}nU(zZHU޻z�� ��i�Ur"�dv�<#�:��c�݋��S�(��Y�̓�M��W�>�{�CD�0#u���͎�N�CD�*v9��k�n��'�ճbk@���c����A����@rv���`6����ٷ����M�Uf��H���q͛ذf����� ��;$�o���]KƒsΊU�>E�S������LBU}�;�6К�ɬ����LR�<�$�ea�j�'�����
*���������:J=�	��߁'<0T���^y�?��� Q�.u�X�Q��ٻd�<����2���w� |T&۞���M�uH$�����ذ|��i���SW:�n��I|x���btz�"�T�l�f-�i�0�2V�&Xο	��D�.���>���g�Rx��5��$4��=(�B.���y�U��Q�����,�)���LB�H����j������%��Đ��b��֧UT�U�Ǉ��U�jTЛ�3y]& m��V"��9Yr�(H�:��^���I�[��BW�B&��.�dF�;�Rގ�n��{ɸ���O��:H�W;y�K�b���<6UE�؞X�]�Id�hG�4߭�*SL�sP�m��]|\�F9=�nb\Xň���s���;��-+�������7CdZ��F�{�0�����k�������yM�3���פ�U�a�-��N�k�%�?���H�ky��ŦO�Oҵ(i���$1%8g�6�+Z0-��kG���^H?_��Q�%p5O\=�᢬�+�'l�A���2�!��ܖ���o6�<�7<	r�Y(ԁ��� Ą}ٳ2�v��)���=i��cR!ߙ�,���GO8l��|���&��R֔�	NZ"�����(@��]I#.�M�u82i��4�����gwL�x���^뫎lah<.B�<�
s�(^t���9��`y�0Kx���Pۙ���=���@�9^��s2��uX!Y�}c�Xw�;�/&e���aW-W��#~H41�iͦc>����v2�t�OhK�����]�eT7�Z���Q�DB%]P�sZ��oYh�b��'�7��N�ϒ��ڝ���ů���o��G{~RKq�	�!�n*
/����(���~��*�!	��>�S���3��J��Ue$�1leyh���Y�	1���΄G�����B��V��l�b�I����e�����&����ę�7��CD��q:�oʑtP�Y�m���D1��\.��=�hk��1sSt���Zt����4���
�� �i�.J��u(+��'�W<`ۓvq��b|�hR�͐����l�P� �ŭ lAT���S���p_�"v}�	�Z��Zx'�	�/�˷�1E��)1���P��d���>������U����	H�LN�q$�s{_�]�N�m܇����p�w��~�s�Ƈ���EX�=3~'�#s��y	�Inl*J��'£q0�Q 1
y:W�� :M '�f��\��y�hġLJ��*���s��!UAq�{�Rj[��� �ȼ>�L�Vfz�`b!%��$��wv*[�n��m���K_�>��{���%�E%%���}���g<c�:�����T����e�a4��r��P
�ӂ"�!��Z�ٕ��ȭ"��V"cA?_�Mw�z=��)IȽ%�,�4�t����g}TF���J.5�������9�	H�OGdK*��K�|��K3!}�#�b�J���ݔa����M�btOvQ_��XS1���(�{��2M������#F?�`O�Aw�H �PI�30+YG�AY.K T��E��yVs���������}�O�D���tD�nLgtN��mY壝��Q���啨�����dy1wh��yh�آ�fPF�b�i�9����'I9a��>照p1�iz���bԼ���/ʕ�ć՛�7����C��QYF�^�|�|E�ύ�I���^�ֽ��B;�6o�5|��z�q7_? �y�9�[/�A�9���#�ӎ��q� ڰ�~�;���#��=�O���v�_&�Z?ָ�br#��?�>k��tv�<�
�x�o4���
!���e����y96����ϐ}�g��Z��y�m&Y�G�O�܄�PA~�ug��D:P^��5�� Y;V�x�����9��6S<o��{��fR�^��cao��P�h6���G�;i�:E�KsUsۄ�c��F�qD�P�ep�|��׶Ɍy���	����rn��o�R��	�"�����U  m��񇾟Әf"���z�p�*Kd�2�H5��0l�yC��*�_��"�u��:��X�N��Y2�L/�����^�{���'���z�]�*��ڑ�Z�Iõ�G�-�MKG�3f����:�HA�D�(���RT�cM۔7���[S��}�;���������3��tl>R疹����F�[l�'���Brb$k�X������i�n���V����@�������a��0{�R]y�s<����1+�q_Ѹ��"9:��,�/u��l|esP������o@h���M*�2��ߊog;�B�z^3��b(�4����(j�7�Sx�ϖ5�R$BUg)T���!6ta�alQ���Rd�딐K���M*�����٘6�qJ��2D��rBҞ
ފ������s��jT�$xG�=�c�o0��η6�kn���4�7'��-K��ӁX� ��0�����Rz�C
 X`�ɣޗ-�d,Jm��Ĳ>[L�xɮ֛O�v�Pk�>�Y��5�	C�6�*��/�	ê
ǩe�I���j��/~��Ü���yc�a�H���v-���1[����g�߬�'����������nƽ3���§_C?P�PB�*s�<�JȲF�3�G�:�o�<���u��rL�FѲ_b�f���}w��3(Ŭ��4U�{z�JtU�T�]L���I>�ĞA�����n������7ņ���V&�� `�w+?��ڋ��Q�%�/#c_I��ܬ�m�8��]�儬�,'�%6��>��/�a����w
o�~*��~�y��毟{)5t��we�0h�z��� �c�]�׹E���H���-�o��Є�&f����#�n��p
�+���B�]Ð����{��H�!L5o��3hJIj�6uU��ԛ��3����(�p�f��y��H�9�bٴ�4]~�T`72��xt���f��+9% %�1��\
qH���4�����+��iy=x�άa|���&�5�)v��1@���R��uIif���f�Ϗ�B�Ҭl��� �B�їɸ:4s0G,di��|�v��-�1��*�<������LE����Nv�E"��oc�;�&B��q��,2�x���,�W�aЏ^�v�{����'��.��,1��v#��[�:hl6g���شν�,��%(�N+�z}��Ǚ��P��+�{2j?��;e�ۼ��&M����d������g��O�f���Yt��_�RX_����`k���8��D�J6|�Ԅ��0n�W�M�\��v�:��k�ӓ�wi�`����#/�*{9�S��� ⛞R�X<E�z� ��W,[�۪]�W1A�y��P���$�z�_0d}c��Nu�"�k�S�9�}) O�@1��W���t��E�����ԺW���]��Yap�Bn��-���)��"�!���g���L?�e�T<��	-_�ؒF�_����y�N$i	���(�Ϳ��]���U�c���S��w-��(c��l�żi�n��$廩����T�����3�C\3�����Xq�G��1��Flb�J6��⹲��`L�&z��OP�yrR7�a<L�*\����9)_V��Ռ�v�N��Љw� CO� �`~�Y����,!���ь�I�P�"�~����N�hcYu���`d{q��V��7��?�z`* ���W����A�B�C����[8���5c��J�n���Hh���~�.� |��+	<M��`.�7~�2$��7��5yE���α���%�Ӧ�(kN���I!�I��7����	�e��K����*c\�8hsa�TiNhi��o��P���ܧ�W��?.����~ֵ��ގZv�u���
<�v?�ֽ54 ���W Օ��-'Z��c�f����`���t"2��?WM)��!�0�C��B�P8Rq���Aә��8	t�[ml����+��0�(?��0T����AcF�*��_h\	��0����@�����ϟ8�
Q!�@4�u�%�� ��������p�\(�by�q��vaLA3.��U ��"5�1������zu��I(([n'Z6��Q���\o��+�{�?��$��}(jta/Q^�-�w�*��`���/6���ذ!z������<����5���ɗ�&��X�-�?��KZF�,tфʁ
 �����g&5!��{Qz��A#՘7Z��Ƚ��1m\��g��w��bOW�W�r��V�3���d=.a�8"�8�Zޖ��LA��ͨO1��˿ݻ��u��&|M�����m�{:��j�� dgoC���UG'�m\x��焇�5��[�^2��F'�sG�@�D���i5���+�`����v��I�dheo������2�La�'t�u8؇]t�H(���]�V�Z:W�D��zi�lu9)k�+��3�'�MWB���l�8Ew�&ݐ�$Hk]��n�����)4[���Qpl��s��/��j�e�+y�C�V����!���Zg�U��<и��[�����Tq��n�k7��~|��׌�t�3�Q�rVF�l�U1�6B���[S��R��~���I�z!�/pha�����j��Q��������]^��G=�2q���Ӵǣ�V%�+)W0�_FC�Tm�t�6%�d�:El���`y���p��X��3#�$�'���q�ޢ�p�7K���k�Ֆ����;�;�3�^U����u���"�J�T�׉����o@eg6���Б�ҩ���J�r��Y���.�\'x�,�r�*��Mm��8K�1
ۏ�;@9BE��`1�ԇ��Φ�܎�0Z̚����Z =i�y�;�_��?ݚ#_�Y���jF#�W�$%��%���(���O��N�L�xU]c����Q��|
<¦�vv ө1�L9:�&Q��\T	���@�n�|���j������ƫt�p,Ź�I�d��� ��	�t���Ȕ^�z��0��0u��-�%Ok�XG�2K����Ē�eX�|��4R(q��dO�������	��.{쒒�������vM���Т�A$����%;�r��&W��VD4@�Ɍ���@,kO=��O�FHQ��	t���;���-f��jQ�2�B<�6E���6�K�i}�����9?/@V	C^��Z_���/�v*m�����[�f����Y�4�����Ѯ聬��]F�*��/���U�m��d��u$�R�::2d%�F�I�[��(!G_���m��/���;�#P�����oM��~K�Qˠ}�ެ�KR����Li����"�=ؤ��y+�A	y)s�ՠ�F��M8�F�V4�l�7=�Xn/=J
L����n@�I>�Σ�����4�Xn�G��	tP�P�P���;p,�@o"w�s�%\5DN��Hi�/��$>�MSf	%���ʰX<��T�/�p Mmk�1^y'h�m���,'H�,��q����зn/�8#��%%��au~�A�;��{�{'9���۹ה�Rr��uo��̹r������Ո�(��\e�i >��p�!�Dp{L�U����TZ*�
m���:֝1"�[�#��Z'�؆s� h����M6/ҋ@��w��o��H���"R�2��X�\�s����x-q5e�
�豉_Ϸ�[Z��������#�*��\�ֻ�n�p����]f|��m�m�3H¬fi��H㛨�^YP�W��`�F9�j$�C1��]űs�Gyb�[(�*���@^O���%������dt+�j�~+!]�����^�&J�a�o�X=s
���F�Y�c��*_2H�8re�2�%8R2� ����)¹�$��˖�G2�f�7 ᄻ�ޚ��*!9H߆�
#We���n�U�Jd	X0���]�~�ο���@v�ܬu�:YYe=w��j� �X-��o��?����'��{�vvK�*j-���QH&�	�cX�g�JC��Is��Б��'}�΂�Z&Џ�T�>RfgQ��o{�=�l'���.��=t��/��@h�u�u��KB:?�X�à�OUq�����b����{Rtnh&:����b�~��+�k0���A�����̽y:;)!��D�5�H��D���!��'}�K3��G;����3[���ۦ���$əb� f�k��$��p���_ d�ttϮ�;��c�F�
/�+��̊SY.S.k�$�&�k�(9<e3+�fi�9�밲d�S*R���>�W+���_��U��+�>T�Ӄi���8�{(XH��������@:�%���Y%���Ϩ�)/�K4��/�%5N�+B��������=L����ʭfSc�Sob���w�d�,a��	���q%<�Jt��N(<�ij'�j�;ǧ�
���>��Vt�[�`��\QN��H��%O��<����Uul�LM^��P-���:c6�X~�B2�n��Gl8�\�S��,�~lD)�gs읞^�. ��I}n�}UT+s�Uzܘa�
ti��"5�trl���>Oe�J5ɂW{�c,��Ȳ��%/)�\�I�x@i���\���^���D�'?0=��#N�ڦ��\˩�h�D+��H+Fj�
���N�{A�~�6�GS;�D�ͼ�t*�j�|�,,&~�H�و���~�3�oy)U}	��TL�h��&�)�;P�*���g��S��Z��p4�լ~lw����ғD��~'}a
h����VD1Y��屮� i�9�
�ޑhN%���]���F�.`����:E�3�6T��꫗\\�̂��s��/�|�5:���C��������*�W��(��V�)r�"<��L�NT(k�I�+P��J� �_�7B(iB�^�m4)��qK3:�$��2��:�Ci�µ	V���3e6�/�p{�iv�����˸'%��um���*�V���&A��Z��wx�F�p�Ǉ�Xhg(dvMn)4hd�C0�l��` {MJ
Y�p�'g�ͦOe	q��88�݊�!�p I���>��k�٨������~S�`�)Α��Q��$U��5���)�!8�~�uZʕ{9R[�)
�ꚞ:�@9���)R��b��Y��R��q�QΏ��.G~[ �فWj�����y`�I7h+�G>���g�黻3��ٸ_:���%��E�L>��;�7v�Z	m=V	'[���!�/�A�6�T�&}-���]�7G��:g��tGEXǙ,k�ǄY�N��P���|4�X�M�va�
VY��x��	t��<�Ք�蔗�ґ�b§ 8d�@�tD��f��W��[��C$e�����5X�Ɨ#	��T��yR؅���	�7f`��q�3��o_�t��g��/������);���b��|�J+��"D��(U�\�� ��}�*]/�;b��V���T�6�l�6r�4�n5�Y�i{�O�=��R(��O{������#En�<OSY����!���.����L��]G3���:��
�I"۶as8W)�<�*4���A�P���W3��|�VÝ�{U�3��ab���Ut͝��7r��oך� ��ڬ�3� ����T�L������c����wXKIk�9����Sg�^֔�k�Bf�`>�H��X�2����|:���Ӹs�k$&� (����Vs�'b��B����$��$��N�K�C7�j+�U%Xl+��E1`���6>Ё$`�����X�f�>b�1��/<g��k�	f�٢y=@�~c��_����,p�I�_a���U�gr@��r�,���M�uת~s�U�ts�o1����N���x�w�h�Y:����T�n��ђ��R��-�o@���t����!��_f� �0�Ɨ�Xdҁ��m��G�n'��8p��w�b>�u0_g]���w�^^��gY��j����7�z�r����Ƣ;P�:RgŜ
�pgw�{��>e_9�(9-)�9�1E�%���`䢌��ǝ	��hqZ�h����<;K ����[)�N�^	��؟u%� x���vAW?�%�$�+cꔩ��2�;sMG������	�ӣ�� ��a��mL��W=5��D��^`.$7��?\�e���0g��z.L����� v�N�d�hHN���<V��y�\�M����M�6R��e:��,�+sz~��܅���w�U��汅��O0���L)1��Xx�E=��iysd~���('���B�Gc�WB�k�� ��^&�%�t���Vq������+a��p��0K��[��
W6�`����{�$�L��C�������u�UL�;>��X,��p8"���Ghy���}!�ʸo��w".\2��V��Ƙ�m��A��}5�c~�>�_e���Gp�Ҍ�t+�!ѶΉ
��Oݷ���y� jΦ{?6�5Ia����N�)'��9RBКj?b�%5啖�����RGw�a3\ݣ@��ay��%I����)��^!^=5�,�n�Ȕ��a� �0�X��=U�u���}��,.�pDSj���!�Mr� �Yde4�'Jo �'�k�� 3[!�<gT�Ѥ>!!���wT�!���d}��4n���Zz�n������E�P���[+މ�2�a=�(���y��dٸS^zd^ɉ���3I�����@M�v��8��2n.j�*��Q>o�Q�n"����m�ZN\J|��E�z��*��TG7�עF��c�xeQ�zR�@��[3s�#I�Ґ��׊�?�
4���Օ%�E2!�����=��C��������n�/A:1�0��q�I&Nm?jנap�,���uY���g$Q�F|r���	�u��@Q@�����4��T�*&7��Q���Xw��%��)GH��M'�ˎ"�و�����^;9���a�ײǶ9��(����+J�W:�ݖs��GG}� ��r����7p�^���V@��&[��8�IU2��>�K6��4	�Nă">=�C��׿��5Z칳��0.u�S?lG�[�Z�l1�{z�k�E����]�2	�%�M�K��9���Ŏ? ��g�n�Dw�,/�|�}�[؀�Kxz;ٲbg�<q���gr%�nSN|�����V�>�F/x6Ĕaٮ�i�,z6}P�{|k�Y��7�R�>�jDBWc�pq����{�ӏ�fO����A�nq�l�0�����Z<�6ٻ
�Y��{�}�FC�cx����d��)h��"��v:)����G�m.�eE�
�G�o^LH��nf���;�ٚJ:B�^�S�B.�qe�č�%��<�w6�����=P:V`��k [s)4������JG9p���L���U�I7A�������;�[�<���І���	��8<���������ɲ�2Z6�CD�l�m�,�S�].�ۀa�:���Vєo�uU���שi��L���� ��k�fĶ���p���A��1�y�' +��G�4L���(���}�!�e[�g�j�� h��>�O�zYb���[�oGDDv�.�����M� `�$3<BJ)���k
bcC�r��=�gӠ�?��A!_�eej_1E����ǈ�i�H"1R��]*E++�U�8�>g;��uD��Gsea�A����W[��� ����D��40h�=�W����n�v`p��=F�=h,N<t��Z��]�u���c�.���҃}�)��*��ŕ����cY�c�h�h�_a;r�`�)!����PJ0� H~K����[���T�u��KH��b%�|X$'"8�{�<U縷Xji�,Z�z P.���H#|LX}�)҃���2sٺvW
����ݭn�!K���5�.WuV-��N�����$��22�����&@�]90M_��J�".����o=腻1��@����7-͔�<)l���b� ��ǧ����g;��x*���{�Ѵ���B�|��{�`q����q�Kg�q͛�4Iز�����n�� c�,��^��Azv��$-����W����Yvn�+�H
ޚ�G��ۇ	A�N�K=/m׻Y/�S���ύ�����XV��4e���-��<����Կ��ꓑ��
��E췪��}�d�S�R���I�x��Z(J����װ�	Kb��-O}�~�`�0=�=��SFjr������<�,�׏�+�\'��Ԁ�iM��ՕR�U5�->-�,�gKi%T}\�_��3����0�<<�	�/����k� -3��7G��Za|!�~b�Y�7"�vIEڭD�8f%�A���?�vUU=Gq��@~VUM+8���ޜ,6|b���~�qn��#�f�l��:�H2�vt��6j�E̻���?�;�U<���m
Q"+Qhax.t1��ǵ�Yz�f��M/sx�l��J�Ӵ�1V;m-�v�n}/��<�?�{vp��ZC�[�eX����%��v������擏���'o�O�ms
j�+Q�v�*���\*x
u�t�1�4=n r{`����Jl�C��*T��~'R���W������� <��5�9�eL��٣Ҥ'L��]XZ,1cI��Y��u��ct��]��-%��&�v�.�e r}�����U�������(���ru��;����$Q\̶�ȗ��-3T0����R}tfX��f�?ۤ^�Z(r�u6� ���G(�
�'֚��ܯ"Y'|`C��[�~���(SЯ�wy������C�=��u�|^�;M�N&Kz�k�
�d0�?�U�RC����AT���WAC}η,����;���O!����J&�C����Ӑu��T��v�{@9%*gVJ�L$c#�y�U�����&�-1��sY,%;�O\O{�� @����fo���#
\�7�û~|y��/T�_�D� 9��s�i��++�/����\"t�h����Hrqf-[�'�k�
�ʔT���V�ف7�+�Ϧ�W�a��͋U��~:J�m�m���NR�3�?]��z�[+�\����0�y|�L�o�S-Djb�.�h��f��H�ت��Tn���3c�\��'k�}��@�
�lIF:��B'�5��*��T��|PF��]�~1x%�q5�g�%k�i��
͑e�
������,Xݐ��|L�s�6�����H,�r9���l+����y��F����	�̐����ڜ�d���#����}��N"(4�������2	ͭJ�r�{U�OƂ���җˏib�d�\��
^��"��A`��W q i1>�c����<�����	p�y3�Φ<	��U�jc�7Œ�o�W
v��-2��j���A-�w����6)�Y�j�N�Q���o͍��Ę,�|I^��ucՆct:�raY�w.�D����U/R�4pՈ[�+���t@�F��q���Lz�c�Pd�����	�k���B�\��-�>�Sk�p ��	`��A������Җ"ٍ�+,�&��7sЉ����#�{6&B���W�@� �����y�hw�'WH'o�Xcv������	F�ɑ���E��~�j�	��WR���FD�3 ��m�jll�ONkIti#^�blCm�b�3�2Zَ	:*�ilƅҒ�ץ't��t�B�����?S���`�H%�Oʕ+��񏛒����D�L_��hl))yJ0B6�Ҍ��V'9�4L�JJQ.��I�V�ٛTZe-4��8��9��p�� �"q����R͍k;{+�&Ҋ�%��#9FS�M������|��{�M���Q�(��D�9�8#�j.g޵~��=��Ǥ(De�+�Kl���X=Yl:���Cx�{�@�Y��X!u�]<n]�9>(����9c>�3_������]b�me7�"�N��$,�~���n�e��ڮ��4�)N;lG����<�����S�`����;�N��Z�!��#.F`��J#䎥O�"��|n���y'�S{��8�5�{)�&�����='$UB����	fE@�ɭ����x�\�����*�z�7a�z/>l��}z}ޓ�]�f������o<L����c�Z:˽�g~������|.?P�@�����<�u4��Na���0�J�+D9(���u&��<-5/�JڤESw�c�o/H��Z��~��y���K��-�;���
��.gc� u���@U���<I��>����s�$wls�YJ잚]u�j�������U�9�lfehr����4JH�SU��&�I�Z�Z\��u\|Yi��H˨���\�i}��U,�:�5�o��s{�8��v�TN�lX+�H�G��@�@5�D'm�z�"��8n����Ж>�g��l�5'�bvj;E�F��p�R��� MŢ/������fC�X�2���h���Ou:����P�ƌkyc[M��@ʑQU�%J��5PO(�u��E;p��w@臀kw ��W���]AzA��K�3�Y�8��i,��	�js'�v���4L��&���S%,@ � �E�H�f���A�#�ך��������x/3L��NG��>�æ��GW��,gN��3~����$PBM�ϻ�� ��� Q��\��~\TD��՟р���m��5f�!z��l���
R�:�gPL�1�*yZy+填w�6��f-b2�7�-�E�wǸ��z��Gվ�Ed���������l�����Ҙ�<�gVI�4K$�	��[{:d��F�U���f�ʸ�@�Ȯ�8b�@��03�i�*���	�5d]��8�h���o!��g�<�Y-�>��y�S�\1�I��������=�]�(���\�r�}�W�	�ׇ�a허^�"m %${E�:Zܬ0�,1/��Pp�Qqq�l��_ ��F�z@yӣB`�Q�@�fr�MQ��x��ά�^u��I-��@��?��~�g�U]� ��]������O1ht�֊$d�+75���o��Nuy����F
�\�MI��V����P��(�Y���d:���7D����;��e-�ͰA���8}`I�2P�x&bk�W�w�A]��/��a����IX��f]͵����f�[Z�n܇(�"�n�j��M!��\�T�Y}`	�ѪD�1�[�a���_i\�&/K4W��0
���1 �쾻f�� �C#%Xh/�Zn*���´��ي�� U)���C�{!c��Od]%����A�:����D��H�?�K`E���ҚQ�wBz}#�]�$�"M�?De���KY�=�m���K��)��bE����Ă8��Q�M�zq��aCڅ}u��P6�/s��9>תh(U��>��e�YY�)������h���?�Ͷ	O���6�;<��h�8��R9M?�@��\�uyf����\����t�:7���QT�5��J�'�K7�r/�ob�\�����.Ԩ�ψ��]��1�,�	� /C���H��������3���)��ꥬ95��ѷ*�;W�w5I+�����Tʣ[2%�g�3�8�t��K�i� l�i#�F��;��#���ơ����_6���nE����]���RcֿBҖT����8>��O�7��]�8(����^+�M��X��>mרɆ�X·�� L����)㛶��Z7�!�4m�ɼ�R�|?�e�^�ҝ��m�1�D����Wg~�%5n���!��|��A�O��������B���fJY���n!�u��a��)yV��޲4wog�������t0&r�i ?�W��稵' ��Y�n"�9���i>i�C����q@�R�3=/�nT5�i���� �c�Q���[�c�*҉R�M�l�}�4GjfG�������w�[ۛ~Yx��ᬺ�P�Z�U�!EGE2>�3��rA|a��we�ؓ��vY2�������'���cذ	�_R?��8�������Dxk���y��\u��6�N푠����}�C���Y�`�����\�
��БT��y��U���NK��[����*I�ϥ��jT	��D޳�1�v�P��Tfq�Ep<�K%H��T�~XI�S��LS��1�/qA%������55���4�R�K�� �y��8�Y�V�S�<�H����~�l������7���^(���o5�����Q���a��Wh `q�`�R�;h�iCg��?��`����\�M�U�lH���o�8*�j�9���bЃ�t���]ԙ^���\�U�N}�a��܏��8L]����ׇm^��^��y�Sx�.�M�}GoQJUtTiW<�9�1������~x��S�d����xWҌ�GYYۉc7�v+c�) �$�J�~�?o�LP���Mt��h��:R��K]�x�R/�w�ZᲪ�\���k�k7��I��4�\$�xC"��<S�3��#�Mq�C��zi�7wa���j�)⢷���Ǆ>[�ǹt�Xo����z-�w��/-��U��qqf�.y�w�Qك��@�Y���`�jG����jCT�GX;���8Q^��&,�d2UKPĩ[1LN�z @��fP(�ORDbg/`���>i�*��Ï;FK���ϑ�٧"���u�dT[�.�n�td9��':z�!$�=`�&]6��(>
����t#��N���/�m�@� ���$UײA�%��"w��BQ2\m��Y�g#����"������M$B�d��Fn�bő"A�d�f�1Mؑ�^9��,���n#��͠K���S��EG�����|��`��t�D��Md�m&�u߄+ �s屈���_(�}d���/�`�C�C�|����yY�{pۄ��	F:���"R���9��6�u�L�f�^~S��#~.)�e�W Ʃ������3?^JӒ� ��|��?Q���qߢ���Q׉�(���~`�k��K���f�aY�ǂ�)/�YM�����0���t�v�$Q�kX����,Oa�0p�3�����v��`]��]�"�FmULOx];��C��8�YE��Ͱ��	ɕh��Z�*��E[��u��JL����P;��.�(��%�6��pm��t�'q�]�E�b(���8�39��CV��\K��'�4��*D���Q����"���&ϐy�����\��8���*j��&$�V�q^ �������9B?Y.[J�%f�E\�����"����(�q)8{x��;�9��ö�+�}f�(o��M�ڒof�J� �\D!Ĝg���m�Ȋ�V�qL{��I�T88�#����]�H�I�&uhI���a�'q�N��t�+0���R���Quiov���|i�P�Z�<��U�z�5n�K��F���|޿z��x�C���|o�p��%�y��MT����'/ZY6�K�Ȫ�۳Uܷ"]�J���[{mM$E�qyq�Gn
Y0�83��/"�J��S7	�q��m�$m*SY�HC��'�|�� 7e
�8�����$���\F�бY�h�J�^�śV�>C��-�BM/�љ�T�FT{Z����yC�Ϊ��eI~�L|�ɹ&E��Z���>�" ��@8̺R���� �s��(��a���/�ia��m���Qwi�{�	'+IڶĢK��v@��=y-�c?6��-���͌��"�fZ��R�<[�>Vm$/W�Qt�d� ���En�(S�5��oD�e��़}"�se9�s5e�W�(52��zr��ͳ�~"]� �xEr����bXk����u%͔��?Z�P��U��Svl��c�E�*�P203���({��/�2^6�_<dig.nT��L�>�h:�L#'�ٲ����^.�B�*�<˔.~�y���m9�!nB|4fq����V'}�����-`2��p �����Z~a%`�n�̚��ʀ���#����JZ,$z	��`$��[}T����x���]�5�L�>od��%B}%�M^/7c�*�eߙn��^B�[���6��ʌJ��o��JN���{���%va�c=�� (��<�Z�['�DƦ�X�[�ۻ��c!*g�+�#5�˅@��A-�t炝��ii ����L�_�ސ�~Z?5�9�ڰ�0���h�8_�{:l����jܮY#����3���T^R�����*9��`ٿp[
�H�w��"��W)9�N�'��i	|Ԣ�_�d�iݒ��Ƹ� ����"UUi���,����;s��k����6�<t|��S��*D`���Q�A�m,@ v�n����>8��|/�&�bX�-�k��bEu�qELH�\����O$h�����^��S�`N�2�a�"�(�H)�^��$������G�m�jmx�Oʗ��
-���,�����iT��R��v�QN!�n�`a�w8H�b�Za�^Z�̵a�H�d��x/&�v����ƨ~4��&����BQ�|��h�HΩ�?y���'�Wьu�X�%'P��*�/t��wAP�k�[���q)(B�Xߑ�?]h�x��e��^�(�vEηF���|T��s���T�v�	�����>�1R��e��}�S����@M-V��qG������Nb���;7�{�>��	1�����͟�m��&Hn/��+�a�����hEp`��SM�2AéVp㡞�;�Hq;;�ٻ�k�I7��]��&�y��%���	����sm���J�5P�E��B̞\�̋E�oi�5v_�����/�!C]7�1+��.	\�"f�vp�i�-7O��P���57�B��7�b���C��_Mf.�L�SP�τ�]���@�߾���G�����W�P���:�p�NdT0@X)����=�e�y�V�bp���/�Џg��(�se�p���eG퉠3jFTDF5�R���i��E��W��/O67
�"T�j��G�&�BD�����p�	�q�5"�s���j���w���x�U��r��d}\*�Z�ɛJ���'��������4����ϩwI����� .�/�4o�֔�i���q��}�\��K+�X��E�-}
��@Cy�<��
6��� ��@��108B�Z�Ѿ�a�������@���9��W��*p3N���[4�*��R��W1p*m$0�M]ۀ�=�i�ֆRv
��D��D�����5Ϲ�n*�D|59Ya{Aj|�6�JjѼ�u���L��Ú�F�)��G/��hoϸ��Xf�Z�`�kN���b��ޮe�7&\r�Z��4`�u��ܩ�)���`�=vKδ��=�uŰ�n	Fg��������?�V����ƪ�Ѫ���͏������>��W� `4�:����2Ñ��G.{#���J~�ae��侟��7&���PPT Pީ��9��<c�07�*5��bn�q���/�ls�{7v���:��9�~wx�sM+�=��b�4����K����
z9��R��[z�β N�*kv�@J ��5z֐ �(r�����F[/�鎦��:�."h�͟���.���r��tGmd�����A�!�Z�RM�����͉�I�o���ne��T����׶�wq�n��GO<?����髯O[�^e��v�e�|ݵ;�>����_�3��>���a�~��v�4���3��Է��,s�!>����Ht�z�������C^��=+.Y��o�=�V~]�H�`��N����蓺4�eOF�<���O�������NzO����!�^p� �=�.WA�\�ek�����T��]J>/(f�������~%U�@+ )�@���^��JO���������[��,�!���n�%�&S�g-��#��2�s)�u�M��ݼU����K8v�HFF���g��.����_5�	�,��` ����FUϨD�a �EN�����y�)�&!�������g'n�0V�����eNͻg���?"W�a����w�(�/ �6���ʉ�%]�uuγ=��۱�卪+�p��w�;�l@هO}K_�]���� k�R���xގ�4=�Dg*�����A�Tv��N���&�Z'�PeZX��{i����QZ214��l{���"ABZ��A��[�)�p�M.�L��uf�0$�slR�V�<j�̗c	֝*�32f*���{ṼJ�@=�-2����Ă.z��7Uo�Yv�@Lת&��s�Jm��gN0=Y$���l�5{���E��Xe��������S���晩�GKD�X/Sca��WQ�f��}����y:�)��kh7�63�z��>o��9��i;�1)�04k�.M MeG�.�H��͍���9Ï��6otTl F��H�Oq[�S�O�� �'�T��mA�9�7�����=�E?�uR�����?^&`�~VB�NR�	���m{�!U�~!��GG��+Y:�Ƭ,si�n/.���/��Nl��&�Y�����J�8%����y�+D�)[v$�B�{�Ւz��fx��sh�����;�_z0T��Q/��r윿�]��vr��WRtEٱU#)?7��浟��e�!��˄-�+ߓk��L߹���M
�F�ܫ�h�td�������sF��f2���c�z�-��v�iCkzD6��_7�}��,�~u>�_%z�
?w�P�̨>�<K�L5��3"����I���:�FU�'�`���,(]�?;'�999pE-W*���l��{���g��\=���;v����!�1q$�{%58����'V��k��kv�;~�mBx6������4�LpJ6]B|����(�X�p�k��^}�-Ūݙ��T�����;wɯx��n���rI/� :5b���4�ET�o���$���}�Z$v�a\�I�LM�K/Z]����U�b�6��N+0F���L� �]�M����7�=��������j��
U?�M�afe�A�ؑ�ۑggtU�u�"n�YA�aJ�W������f��G���`�H�e���\���jd����z)gǕ<'	đ�1��Ed�|f^z}�c�?�eiwjZ.kn|f>��®O�e��������(u���«�~'^��#"t���6�l����֬��]�,M����Qv����ȼJ[L��:��	��y�'y�����,�Ыf�XU�}�3��$ ��K)8�O�Ω�;-q#^�\�v5��&����'���m`W$��fӸ���+�@e{t���U�j#�����j���f 0�>]ZUY�*`A�^ް���1bao����/T�s簠V��p�טPmO��ϕd�|+�6@��^��\�N�E�%���Ml�Z�mޠE�<������
ݯ�ۓJ�������C.w��Niၕn��^Vy�N75E�ѲKq(���y�NR��nO�v���>e�.t�������r{'��F(���ʥb9YZQ�F[r�2[WFxFm��S:���n�N�o��1����5��|hb~��O��jצo��QJ�y4�wj��;CVF\bf``ly"�0BY�:�w̶�D�I��]���ۼD����o)��b�ϓ��`|U0;+�w�#��tHq^MPh�H�3, �1�����hA����>�%ć����~��	l/-�	_�ō��h8,�L�jKt_���&MQ���H���# �.4+2�ĔE	���_ۉ��ж�f��������O}5���_T|X���+uS�q|�Sr>��9	%c~~и[w�*s�[���ˈ�3��W��D�IȉK�Qg"GA!��!�\���c9����o��q)ї��z"��5<��6L�Zm�!���"�Yj�5w��[��V`\��lδV�?<�E��Wǥ4v@��ǩA��*=�����Oc����Xk�{Y<Q>fȫy�P�C�6F���"5�;���D��5ry��b6>*<�O�tF��/�;��'%'��m���q�{�-�����0 ]aZ.<�g8t	*w���H28��R��{�s����0��%I�ل)Y8K͹sJ����m��v��٬�-��K���6��N� yMO�C0��O��lW'^�K�|Fȣ�`�V�~���-�=H�����钝Rr��:��	�g]�t��R-MH0t��b@p�lBJQ��G�'37{��i�-<w�i�J�&Q�*���潊��<7票��h8�7�<�'a/��ZV�<e���0]%���J[*f^[��8���+$NYMY�ti�B!����P�o�/9wN��Ze��J7�+��2���R��ލ��f�5�o[zTC��Κ��a�
�����!YIe��~���yi�׻f�qJ����!�F�����T��7���c�B�4Z��_{���������x�ʹ�P38����9df|h�d�g����ګLW��c����O�Kq{7öжS���Va+�i&uW|�2��?[k�s|���G�����1�'�MP����1�0>��#k�  �u�h�%��"pU>�l�c a��R�X�������`�7����	V��:P�[�C�(I6O��,U�W�
��3̀4��u����1�����'X�Y�� kE�|p��0f�q��l���[��M;Tͽ�U8v2����W�~��-� �}ZS1�ly6�2�Y�|J�`�z����ŨQ�wI:=2�㛗V�:������.$�����"՟�X.5�څZ�W����ѓ~ijP�{�ڤ��K�18�qv�h��oO<_�eϝ[e՞\���N�Sl���A�8z�3H
�"�R�-�ۻ{�� *w�J�U�"�d�8\7�������&��׼�i��V61�W 3*v����$�c=\����݉�FԬ��^>�i1����w&�-*�˂nVwC�!G,_��C�@:8U��9��|�+�x���
 z�ر�:��i6YAT�?�����#|"�s]zl�Xd��R:�V�S��-;]�0�6E��9�ا�L-]��7�A��]5Ko������E�d����f*q`�92�/~��b�Y�p��8!*yS���,穞��h�Bu8� Q��1鎄�e"u[�� ���a���c���gz���Vt�O+�8;��1Ю��i��f#'�HPg�៶r��`�+�Y���-�)D���E?���4�&����˻����O���B*���"`^���,��,EA����8�E-�s[*�6���#�S#}�M�٠灥��ˢ��� "�`��<��9`����b|�]�;W�lY9W��kݑ+Lb�����@�kD���0�itH�-k�e��}��T]q��l>��h�K%ۯ[��HD�<�Уr�jl��_�\:I%O�$��6�{j5�������KyySڻ�"S۔�%���!��N-D �yu�^�80���5~�˿�N�d���d~������W��8s�T�d�k.�A��J�4VC��N/�6?�f�U*�ku�g	�H�d±� 7a�ȸ5��xξ	ao���m�B]�:�W�w�v���m����;�p�m��bt{�^���H Bd\�X�UM��A��?��DX����B�8�(ɼ"���{;���+�4��d�էJk#:�W�u�(�n����U�ۂR8e���L�|��5����a�X5|d��t{M9�wd�#�� X�gZ�*z��l,����z^�£�sŷ:j���VR��vj�]�%0����=��Q6�l��L�c���p��ļ����t�u@n��X�|%~���Fc���z-o���b_�i�:0  |G��bѕ�Te��Nbm6�A����vf������^z፨�"j��z4��m�֠��R!�/��<�����'���E��϶�<&������8H��G'�#��@A��R��|��k��,�;������L�r-�f/-=m��FM]JvQp!�n_�6��FB���	�Gxa�?=��*��.�n�A�u�B��ܰ����"�K��B���"�Ԣ$ ���ѕ$'Զ���K�hy�j)�K�+hɩL\�G֣l���Zl�!Y�H�����w��J�@Q+^��J��C;gɩ1ҳ|k�]yËm/l�@3�Μ퍛xW��&bz��N�m�/_�seh�n����a�t�&�y���<�)�����1@c�/�ъǠ���i�k�Y��c~�#B9���ǥBvh�-�m���`S�RF��c� �+��)+Ժ���oI�!�U{�2R�ڶڲ����(7/���t��Ԥ����@@�X#	ş05xBs�/ܐ����-l1�v�- :�O�p��B%	��`xb�8�X&��]�p#ማC�?Ӌ�wb�A���\����o��r ck�dg���8��q�\V�G����0�?��SX�n�Y1�݌���#�
L���Nz��2|(W�����r�Zz�MI�@�>���f�9r<��r��y�0}ꛒj�����O�����3���=+1}a��6���
��f��|-.�b����Qb[s;�ݟ�'/+2L��m/Nͯ75ϦG�;I�u�=I K&y�V��M��{F�i�C\�d�����󉘴g�u�� �o�l
�:�����#+�
��W�V�{�Oc��.��+l�"Y�/�4�ʅKxȲ��	��hp�<k��u���ʅ���-#O�&�h�sX��H��s�����Ϋ��W.��"qM�� �5=mϠ��g�?Q�������?�Q��&<4Ѿ�XI��gŗ�M"㴲���I.���6�VwK-0&A��'x߾��B���	�K&��l�-����O-Q�d�=,�m��6phH>��~Fu�M;?��\ Cߪ�d��-��}j�ĺ��X�c��J-��ʼa�Q���V�g��Ѥl�%������ԑ@�"����$h�X� N�o%t�6n���^��nQ�rV��:9�F���Ś8U����d�օ��#�f +0���я�V��J��(��!봯#�E3�!A9���B䷐�ڕ֦'T��<�켘�\)<����,zWQ�m�.8�3�q�ר��}�1���k�J�x��E��q��_R+��U��lTS���'��%�i>�����j0���jy����E�4\�����%�@3 ؉�s ��s�6c�����*�������)X�F��}�A����xLq�'b�a�e�V/�]i� h!S�P��[Nx�X;M����d@�ڐ+}K�a���u��
��#�8�Ӛ���5u�g���;�k��б��>�Xp�}A����"�>;mJ`��8,O;f���������
M��ר?x�Unlꔃ<���ouDAq��nX����؋o��:}�-�X
���N�WDK���\ƞ�bl&���8�ۭ^�!d��6Pp�w۰:�Ѐ
������L��k|.8kj� ���|�ƒڮ5�ג�Ծ�8���&�"A�8�p��N�b�P�e�M���Nz�x-�~�*;�oza(��T�%�<����|ܠ��TvNEar�ZVv��6b�3���Fu���%L>�.a����n���6�����H�=BT��)�o;����j�4~qc��ӛ|���N��!`�c�ðO����P�<�-��+�x��$�Ɣ���Ql���=`H�rzg�H��jZ�iD�,G�m��C�ծf���7ݣ�«��:K�%�~/�[��W9��$�pժ���=y��ж���f�2����n%Ff�Ά�d6���J�� a���Q/+ �|�dB�j�+���@�_,�(Ѽ�~�.��T��녅n_E?H*Њ�ֽF�e#����o$�Xd�l���T�n]�]Q�2"=�}-�1I���w��&�wB�ϔ߾�7��}�>�k$�n���_��#,�l��"�xk9�9jy�������#;x�aWp#ޤ�Gp���̅�r��9F�*���!BI���e�I�dP�"�)�� ̛K�� �|�>j�F��^aX%M�s4�6�/���M�x��;]��etٮ��-ЕSc���V"9"e((FX���غVVt8o�nw"��j���#��o~p��tnP���"[0zD�,J@_�|�I�%
ՀYE�~@BD�=���+�r����˥�D�h�����J��h��� ��0\�doN�m�x�Y���˂ء�C�-9���1v$�C�S��m�1$���j����񉞵��Gw]3_�fHq�Eyi�-�n5we�)缀.��ʗ�f7&������L80���*�W���P�¨Ѧ��gǞ_�����'7pҿ���Q�����F4uE@��������}CThnT���Ew�0�H��?�hԲ�01�v(ot���L�/�X�|����#!���y�e��+�����aB�[��-���Yg���D�+�G��N[�\7�J\aW����u�yD92}�.���)1Ѓ���i��ۅ�)LZ դO��ok�$x�q˃��u/(��/Z2�>����'�C ���/�,���SZ�EP��p�4�Y���b�%AY|ղ��쓶E�sV6O�O�8��h-ݣ�{��*���	���]sc[v�2�{��ܞJ)���pf��aRr���QZ�>�s�U��T
��)��$��b�?%odI���7c������j�Z���%M��1p˭�L����
�a�k�
��Lý���i�c�t�o�/��dlJ��<I�D�J�h���B�e�Q\/�ↀ�����c�VR'/D�
-����}e�}�-C�PR Rv���� ��D��{
۫m���Πj��:óp��97�OΈC����᛽DA���W;'�-F,'W�K�Фޓ�9�=�c�Ir2���\�������?�����4�*O����'��֍j7�g"��f��W=m�����l��	��B�)��!�XR�1�#.sqL@�+�]�RK=sA]K�&��DM�M&�`|�ް�w�\�׺.ѝ��u0��I��	T_y�&��c�
���,��n�F�3��))_���cK뿈�'�>��:��`Wݱ*Hw�(׬�����ʽ*�U'3l<��m?��뚽e�i�4f��h:�5��0OVSw!q[}&%7�P�u'ar"S�%�����Nt�j �/C�Ƀ�.��e�px3p��o��m�ʜ�����9{�����H��m'��1[���	d�S�P+n>�N��<A�,1�X>�x����O�X5��I��4��r.�w;�0�nLV��)�U��3��n�[��"](��)�ں��	R�5��`���
r@�ټ��2�ϣ��EzyuT~]�������`-������^�5�p�l��XF�Ʃ�M��2������!H��U?<��N�$B����a�^��u�%ڢySnS���O�6-H������
����i�%W���;��q����g��IԽN��a�2�IJQ�g2d�h��]�����Sz�`��XݣU6�h�ҶO*đNK+1Q4��|���<C�r�8��	���D�:ɺ���i56HA�, �M	�^�p}�>�Y6�=2�>��~<)���ـ��n�6X��o�����
��<��$"��r�^�P	��ūd��N/��X��V���9c��I89Y�hw�H>�y"ſj��:���08}��7��~�x�(dә�ٱpW^�7a��-�[�=��!y���@;��i��+-/2�=�K�����
g_*�6�(f�M&�<.	K�B�;<��++[�`_F��kI(���s�A��� ��½B�Xo�@�f[z���=���Y������Z"Q~�M����}��US'qg�v.�E	(i3�3JaD��R��_?e9���У�gP4jq���ӒEs���/��/Y�P	?����wqOľ�+�V��)��G��G�0����f���:"q]�BwK����S�9���Ђ���n:/�0h2���zz���5No_��$�##B��\*��� �Ȃ�N�0�}!&q������j�u�t ��b�E�c��YH���B�^���P�d�Z��Yn7ط����Ւ�'�9��{�m��3�ց]������k��w���X{���R��>	�����4īLw���t�L9 ���K���N7It�I|e=�v�i͌��il	��(�J���+��6 �����<4*e6)"����f�xb�|�+%���Ȁl�rw�c�RbH8l�)r����[\"�[مj7��6���;��{�#x��E
@�W�ۉ� <�t��-�׶ܵ�m�ɐ@��|��x�7�4���N@���
�#�[bLlE��
"��U��5@ٱR�a�
U�6ݲ���]���O�Q��=��};G�?J�s�P����������2��P�&��L�P�e��W0~��c���q�T*�Q������EGd������x���S�� ��E����t��bh�z�,��fs�a<sm�Di��������L.�R��In�:�YSmJ�:=�e尖;��|�,|�G��,4��a>�_ܟ� �dwOK�K�]�uu�a�̜<����2v��$L%���r} ���;6V�fm�E^"0�8H�Qcʏ�5�NȻ��@�{zOH8�������'g�~!>O�_�s�t��%)�P� �V[F��[�昤�yX���V�H��L�U��Y� t�2Q�����!e�o�	Tz�}L&�݀^w�[Q;�'b`;�~�sM$�MiB��4��
��_#�p �f+N�W�/����0��%!q�/-Lu��Z���z@^_�㍺���PQ�8�y&�,��T䲶|3��E�L�^�
�iŏ�S�BT��/�k�� ��M�j�|8�\��=����TUܞ�d�ܺ���A+�ACaa�=5�紑ĥ�����T��Y��"�S�;��aP�F�]�,Z0s�����5)S�r"a���JC�z�<�/�n��ǧ\��2�v���a �LOMIV���=#Q��6�a�S��fj�1�j��"�O�ՀEaty��Ǿޒ���r�����AO(����A$F��j��Y4�=[��\5b"���$gB�D��LBI�~D����<��0�6F\�K���b�f�����Z��=6	�;'��{��tC���l0���B��esm�O�)�&���Yٟ%�c����Pn�[��;-�]���G,���H�L�Ӻ�ՠ+�Xm �=F�r]Wc���H���F�΀7�|[7kҀ¾)��׫z
�'��&�HC�{��Ń&*Y��J@a5y�q������G����)q�����;�z9��T�'SLe��b��	�ޕaE��t��TuY*��� ��]�莢_�a������z�I�������B�B%��Uȩܿj�]��o���6�wH���V��(��:�Sz�AG��ŗEZ�(a�E���c���=�*�䒒
�~p�c^�y�ߖ�▭<:�>#��C�����S����kGCI�r�o�e�g�cM[�ܵ�xg�w@�F$l,��4V!784	�I; �cM	>%��2�:�����~ZH�<OPFy��XW�@qJ��iyFEG�~B;�젾�IAңu
�ӓ��M�%�ufϨ��_NT�����XO��B�g�^<8�S��?�����0u�5��aQbɵ倒�6{�`ZLҹ+�"�d��a;�M����c<���%�p�f��?�!�`H����C�K�𣔥^%�O���һ_}?���`�X:�g��h�@6�
�o�Ylui�%k�V|��0��)L���7Gp$�uk�
Cm��P|�V\P���L��a��e3 P�8|����C�����@�h8�i!�ͱ�P����������5�U,�TWeg-�c��sJ]D��\���l.��ݑ��o�O���BkA�`N�!�������c��q��q@_���S�H��^���~�ai�B~�B�M���w�lmd+\ ;�b�q@�>���#�M�̞ �'o�f9���i���s������4����G�kZ"����D����v��е���ib��+w�RX����LGq�8C�M/9T3��i����H5f� �{lK�&�څ2=;���NkR|�uŋVV)��Ȯ7f�z8���}{��Tƥ}@%�Pt���s���4p��R��g��)!z�}��b#��� U��C7���A�V�HA�u���w%C�O�2A͢��ܴ<ZAV11LA,�mS�q�@�Ϗ��ym��^i�=�L�﹃J��������bL���IX���g4�,�|�C�-W`kX��fj��X���a�8Ty_�H���-��0	#<�<�k��_MU�TORے�S�ˎ~���Ÿ�k���+�~s&���G%��7q�l�@Y���wr>7G�we<�� '����~��L�g�����5� �m��p.��W5;��>!^D��#ItB���jH�1n��.��xφ�G���t;ڨ���n��L�+
���}v"	Up�w��׳&S�����}@*�_���jWh@��F��,&w��8fg$�*��T��o��"���ǘ����y�a�Th��n������uJt�Τ�¤F��r���$X���.(�Y�MA�,9*���Z�����[f�P(���j1E���zm�R�2c�P�k�E|��ᆏxO�<ׅV�V M����B��+��y�REqD����,��L��^�Qg�KQ���#�͉��{F��J�v#@=���.[����0n�v�%�jƑ��;����������,�(�&!OY44�RQK}�2��j�)�O=S@�U
�B�.�@��V̻!��F�(�C�$�i��S�G�[J^��t���K�k�N���kF��D�o<����PkM5�v?R@��fb`��lQ��\�jq�ы�ٯ�����Ǜ�k���.�#y��ml����9[���ᦏE����������j�q����i���D����벷�9; E�k����\��qg���vO�gO������ 46C���j`�� Q����������fը�1�,���j���I�̰�(o\ڼ$�qFz��}�ʵ�����������,�T�_��#o5���B.�Z�Y�\ņ���&]�MOs{��n�G'NӍ�D�ʛ� ͭn-�V�y4�aZt��x���N;|�s5}!��	�eӉ>��d�l��B�V�e>2Jj��D���)��:�a�͹�L�*����*�x��D�*iGo]��*S1$��2Z��gmiu�A.!R,y?�uҐ[#�dO�^�G���%"�d�#����Щ�� �8t2����Z���l�Gxd�"~|�/F�z�Y8����M{��Ĵ�F����1�1{S_70��	؍&p��2u,Ͱclf�F�bi��_�ֶ��HHuSɌ�kð��JJE��|��Yc7���?���}�hF\�v�*p��gU,}xy�~d�ם�ݽ��*��I��9��ڲ;5a�7B��D��Ǟ��0��<���Qgi#��dB6)v.x��B���7��'��OBt���P�����~z�ϕ��G����Uq���IŪ	:SAHA�4�ѻҙ�:`p~����D�$���<�/-YQ
cE�]_&��`�H^S~-]tJ�UQs�d�f��ӓ�G_h�O1����σ�M��=���' ��.dC���u8WY�
��������Tɤ���Μ��{��V���.էҏ!ͯY�Ło":>�5�ƍծ1��!'��ƱY����&�ae
��Ab!D8;�XzG��CΧ�$�BC.�_,w/p�m�%L����f}���Dc�5q�='��P2  ��̉R�ŕ���k�R�P�잝D�܊=K�I+H||u�8Cuś\�?�j�J�n�B	�@��Z*�̢�}�}��k�|�f�d&��%��G�ܛ���:��G����h��}��j��Erg�u9D�>O?��jL�>뒽@V��r��E�n2	���|�.�H��d�?��.+M^�P1�)O�5!S�t�)�7�:hO��A�4,2e +���{	F��\���*R=�����{CX�[S	b��S�9ѷF�a���XvᰃuҝE־J��F+���S�	Gђ�=�	գ'�$��uR����yuS�Bz�w�b�6W��LYftU����Ub�l��91�9�@�0����l9�����3��r;�_Og���Mv�7�`B��^4 ����Q,~���3t�?��<�����9�}�`�tk�<~�b��L=���o�>w�Q�\ѝ, ��=㫑�}�:���cj�Pޘ��c�Z2��h�������T��A%������c�!�U�_'i��æ�m��EɎ.�ާC�M�?w_D�`"�km��0��%��L�e*�S)ԅ�TD��@��N�22�+���6<����8ߎ5\X�4�����>�<�, �|A�1=	+#��ԌxQg,���̲��:��0�I`aVP�*Q���[
{}n^`�+=|(�{�� >�sw����(#xI����(+g/-�@�`
ĺhP'<�	��t�C�`3�%��w���}6�D���D���2?���捏� �8=�i1�+�Y�KO��5ݔD�|�莧��R�����M�y�K&W�I��q/��A�~�9�d'G������/�u��xKόp7A3���=�vl���,�T��W�hG4�k:�N
WkZ�<�́�R��a��ŰXp�v�<�NP���a�FSAKu��/�ק��hY�IΛj��)܋|�s�𽐂[}�	������3�����Ɔ"V^H�r~L�t� /ң;y=tnR�<žL�SMIl)����Y�\�r�K{��L'��س��%'h�G�?�̞�S��@-X?x��{,8mEk�����F��r�ܘjF�|�;��UYP�M��K6��\eU�=?�{��^�;f[�@U9l]O`?;�	+86!���o�^�s�
/+zo�d0I��}+����Ak�m��b()�BrY�`Hn�ݎ�2�ؒ��Xɫ�ޕ��@����Wp�jl���t�I>��ee�<v\����_�I�\X����� �",.��X(�Ǐk���|���P�a�A����":��9�5yv�ji9(��#ˬ�Q�-��Un)e��6�+idd_�M� Wɉ�O��jڮ	�d*�]�NY�K��0��C�ހ�*#3�"�P��a�KQ��~��f<=|�>؎��)�@�}���_߾>_	.SŤ���obQ^��zaU��-�fB�/Y�q9�`7�N2hr�}�^��p,�64T�fj�k|���%��,?L�'�:� �Yk?U� 3_�Qɏ�R5��>ˎޔ^�mĨ���� Ep]��'�����k�u��3d���?`�`Ef2�[�}C���N]�q*�S�m9,xp�
�n��˕�/��f�"�����*j�)��[fx'�k;��2#o.'
��~�ֲ��@<l��$�lU2�Y,����*o�I9�>l�^�2�<���GQ�8��iew��i�"'?�<2E���ǃ���Г��F�u�}��b����<@�{��ŲJ�l����w�8mx�E^�$y��L���2�À|K7��y4Ѯ����.�U$��M�����\��qu�f�s���hO����˄��'��0-�"��у�>>�Ѥ�}��R�n0D��ώ4�P[���bPT�T�tW����iB�(I�r�������H2�Z�'E��Vy�S>Fw�Y��'8����UYL}�Q6.^'d���ԡ�¨���B{�m5�T~N���TJB��V|��5�X�c����5��lǳ��%\�������P6�]&��:�ZG�U��g���S��]���^6H�ND<��9�O8m��Cj����
�<�^�N�	��7ǅ� '����{H�}��N�ψ$*nmr�HY�?(k��Z�U���M)˨N�i��c-�+W�/td;v�-����Եs �K�N¢�%+�Q���q��aru�W�$L��h�4���u)2�r�ڏa46��1�ῢ�Y��E������&�{��3��!��{�WZ���E�\�%C
'����J����G�:����&��&��ԧ����nF��q&#nE\��2��sjĘ��r��N��5v>t�I^e��	&:����V�:.�ɩ�������z�].P]�7G2@b8K��
x�[XD��Xq���Э!Z�\~�k����d#��#p�	�y����WP�0���w��;Є�1��|{�bG{3^AI�����ϪdR��0k%�P��1��xD�O�T����i�X�q�i�h���6! Z���ߵ32f���@�̥����>� ������39��e��^ɝ:@��l��
�˳"�I�l�P��� iY�^&� ���|���Jl����~�J�O�1P�3�� -��i�c�Z�j����Q����+]Tl����ᖪ�W��!B�Jc����Hu�z����<�$��T��l١�ǁ� qy��3O٤��x�O�]���	3��Z:�o��I�NdQ���d���6[�U7+�RRh]�,�Mcv�� +���u.��8����Ⱥ�b7����8�/���Id�`Q]���p��(���t�KA+NIB�<����92s"��H�ϓf�.L;<�$^��PM���iS�ᶍM�c�b�gz��F(t��$��fn�I��L={w`�xC(X~�Ӫ��}>���m^V�ucG��J�j��D�:G���h�%�Y�#����|����]���V�:��pN�6�2$B�^YB����|���Kc<�i�����Vi`֠u�|Yջ'����B�"���P$�{�t���ett޽�C�h)Ziм�{���\b�d�|�iլ1����O?�ݥ�-]��t�p�k]��7F�%v��tA<���;Ǎ\v,�%�(�KLe(�
��DB�T]�T�Q�97��07U�"���
���i|<H���y��@KA�N�c��߯������Z�ӣ_��&ƾuC���〆��0�pN�/c��0�{�O�]�x�]h��^��1�*U2��?��H�N���W-�u3q��5ؚ��~Ej����ǃ��Vn���v����;�����570G<�� ҆F����>��	G�ȶ�~)f1P�[�.�S�)�E-^MJ@Z�b���S5��=�]X`�h���v�,�*�xp8�3�@��4-9�C��]AȤ��4[#�;!f�����y���	�v#u�#tE��=��N��ĉ`����:ֿ���Pj��r�]_C�.����m������fa-���$X@�q},Ch�@W[���*�uJ8�m�/��H8@
��w�H� �FWT@�H�j�OF�g;DǍ2��C%[`�G���μ6�ъ糖��[�����>̮��xj<5WO��aFK0��:墮��,oΊ��yصGD
�<P,��69�BF��w�ڭ�C�wYR͏9�f�ϻ ���wi�bm��:-�ifŸj�S��B�,Zw�w]��m��I�깙��1rK�$�"�M���؎��X�:`X�C�k+�3�A�2�R�LcQ��3��H`�z��Z(۪����w���FB���?��Xp���zߠ��ݴ����aKWţ!ųm\4>p�b�Ȅh
���P��~�VRkb�2��I�������SK��x�Q�}q�Bd�/����}ba�.����YU]��W�Ad���t_}� ���	l�*]#�}R�~��2��J$C@��@���bl�I��SQ8o�bq���r�8_r�Q'�{r��<����Pʙ�p����������!b`?7b8�Ln����O���DdZn��OR�=��[dK!���dkϜ���哇y�Q�Ü�{��t���$��TT(H$�}��>$��Qs�WW[pƷ F�Y�V[��$���6��dՄ!h�����p�tkg_���-�Q���vnrtYk���Wj(~����GMS�S�'G�1���sǐ���vYg+(Qu(t1���W�m�)��w�8�Z4ph(��?�͙��^s�3�c�y�����Q���N;��T2O}�|_����v���^�� �?f�(�:=���o�����kR��A��J�g��#�������d��}*��&�0jӼ0�0ER��߲������n�͋�l�y
�u��b�`���؟t����E�s����0��<�5��_�e��^�%��Ml����.d^�vNi�'Q�͆/2�F�*äA�.���"w�e��񺮧L��r�N��w��n��7�ҔYh��&I��['S|y�h�w/�{����{�@?	�����-���/�%���ln�s���}��C:S��ߋ�}�$@+����`f����?|K��_o~�t�җ�16*��Y�=~�!N�堣J>`�{��w�>~���m{�R�0���T莢�M�h�� J�q%�4�������N~�16p�wdh�x�j������P���}�᣻y$�FO^��k��v� ���lq_��B��u�\�{���D�R�4'K��Y]ܙ!��^_$�m�u.g>��iá ���I�������/�����h��L����SW���Ȑ-d��H�-��P>�	\���Aue��c໐)����7��r�U�\�f�I���&6B�:��I�S]�X}3з��G���/��ق�௷�a�h8S�E`����[cM�/����X�2Dә}���ᒁ$bQ�KRx+�w5sV4�ŅLAy�0�~^,\(��K'�@�'J����g��t�w��Ī�ow�^Ӌ}3ґc�x+���适��T3��r_}V��j �ݩ��`�Q}�mf�� Jx���=D�G��:J�5�k���~�I�K7�R�X^�����B������	'37�}���b{�2	���o~踆�S[�f�(h��V0�Z���ԊEQ/Bn��]���*�z����u�wY���!��>�T��8�vp���,c�!������%��EiH���*W
��f�
�t�]}~�T�����jI2�.�������-rA2\��-mZ0v�B�8�hҧ.�]�������~�U�>e&@�qh������Z�"Y����с���&�w#쒏�E�	� B�A5��V����+ӆf��{�c"(�\j�Aa��H)��t\�5����c�	����H X�F̀W����O��q�j��w��Q�*�n>�]����6u�������}�ab�!'�=)���\fp"[>��/�s�瞂�z�u���C�ԩ����c�z��������X*��� Zf���m�S��5G�����7��.|_>��2��a.�ۜ�񱼑6Q`;�c�v���#��{��ׯ�� ܸF���I�=@b-^5�k�r7��E�~
�1���-�VC��k�ȏX5��ǯ����W�9�T2���M���!u�=�����e�txp}�dK��y�R�-��^1���~�싊�"�	����m)��|r�|�i ���)`����85a{����?r�V��0�~�5�`����:�^K�5�°lT��
�|�f��=�a
��J�� {� ��ȍ}�-A�zc�	�&bI~b��S���&�ل�!u����+��JR�����~��7l�D#%q|���}P����2) x�u��uS�e�Un��Ky@F�ۧ�
*()�m�[H����� ���D�-�����Z^.���l�*(
$��r����ع�ک��E-�y��Z�ȶ�I���L妗��7Q�	��g4���Tɯ�Ev�n�r�<���Ǿ@��~w5���l��ݠDed��n��B���+?���P���7���������b�?��<�*��`��vj� ��1���q�3P��6��g���@�P��m����
Q�:J�%q�����Eg�|���M&c/<��[s�����턞�/�4��o��������������yo��bXP��'Y����*>���q���H�����a��!tQ��`H��f�qcR���5xΒ,N�8�C0��ZM�������lP�����M6���]lͥJm[҇���t�|R����)�|?���`�zxk��.�,�,�A%�bt�o��+hL�;�ϸ��m]�]��agN�7Tȋ:jN�T �{�쌨!j'�IS֬G�-!��J��C�	t�T �R�	{աë��s���L���{�z�p���U�t�fs��_u��[)�h�Ol�ן�bT�_�,',�L��W�m�E�F()D�Fϭ��<�K�:.�Ĉ?eڂ��Eٷd�%#F��M�D�YB|���b%Y-9�ӇqN:��I�͞"�y<ۮ7"tǆf�����x�U0qo�4��K�����O%�[��J�� !�)�$�e�X���7\�q�̊��A���kY�&Rؽ�`u(9����7�,|Vs9M4��V'h�+(&��3Q��C����3'e}� ��ʖϑ��j�{1���Am*p��5�]2TAz�FR:O|u�f)��D{B�~X�d�,�_p;�;���}|�X�K#��f�U�"�6��7X�X$ybrN(0uccC�}w��6��S9Y���S�bJ����Yh:�bͷ�3͊��������c�#��b���I�[�9���l����G9|�F@�߻%���t�]��r�Q�I��_5�.Y�Ó_u�%KL �u�c��n�	=�(K8���d�ܧV��ul�L0��sY�����H�A��ZA�~�� �ӂ�*d�j�F]{QX�����DeN�խDjk�\��V�K����>�������[r��������h@���,��Φ_\�	���X	H����
JJ���.�U�Dd��ԟî�,	��3+���\� W)����-�W��F�v�ͽ��v� �)X�W#X ��"�h����OܶZO�|�>[f�e�F�Q��f��'�Ѻpf��x\d�d��#l�T�a��~ʦ+�?��ƾB�����@W��
d4h���G`��� ��^�h�Z���R�3���."� F����!I"{�
�D�o⩈�����#�2SFl�����In����2`C���%�Oe�d���A�ʚ��X�vh/������KD�n�s�҉���B��
u٢J:���D)��*��4urW���ᔖV��S����o�'[�����n�M��c�1ݫ��=����m@(m�49�Bǁ�$�SJRn�P5���lu����$j��զW���T���*��O��,���>|�@4Is'�N
d�K�Js���X��V�}��~F]��#Ӈl��xxD�dPX��T{��(�jH�j���ΰ�U�����e�e����B	��+��N���%qN� ����h��7?��=�d�H̽���'����Gq}/?%�I<�10��I�4�|�����qС�;�y��^�\��ݎ'��t<SΑь@S��;�!<S�E�F��d>*O\<�_����� e�>k2�E��t
c9 MRc�d߹�$u�%�P�$�2~�������M�`*����� �i�[s�rm�#63��;jF�T\��g*�	&��wQ�^�-{�0�j�[��AU���O4E�l���L�"g�����T��G؛��U�ګ�߱�,.V;�����6p;G�P��r��n�-k���B��ߗ�L�\�U������W��Yڔ්�P�y��[6D#T!V~X�l��UNֱ�M�iḻP�@�}I9U�%�Wh	�E�y�1L Ɨg�x�qcԵо3=H��O	\4��k�e������Q�uܛK%u{�/T,8n�%ZF�7𩆍���i�sQ�}b����B�(�$�<OO�C������g�Q�	=	������]�\�+�I��ճ�{�� �e ,mfA�kfS��x ����$�c��Q�b㸚n���ܿ�x�{3,	zˉ��vpّ���*0�ZK�ә�c��Te������x[����c�]���z
��{�:��Q�h���˱7I�����8m�¬ �{ҧ�S"���	�6b([�0]2�ku����_��)I�����׫�r����h�1p�d�J���a���LE�8N`&)b�s�-k��GE���m~M�ü΅xx@M�"L�:T@թɯV�7\�4�tD݌�z���q\L��6]/ed�*+ŝ��w�Wئ~�3�3A?�1�����h�h՗�Ht�f��ç��$b�5��AU�͓ �1�����ؚ��{�W��&��,uƂg�t.���Z��k��F�*��x�u1*�C�����OɎ��]8���M��:��oߋ.i�dKx�8��-v��
�����%~B�6	+�ʠ�%�5���ٳ�"�"��{��'\�=����!舥4D�	�8��l�z� &��dDe�J�6E7��ρ����s
�~|)�C-l�z�Q�	��P{��������\�h�����{���P�CI�IĮj����?Qw9n
���r�3��B�ℎ)R�6/G����h{ߐz�ܸ�S1�7�VkյSS���2t���U{�;�xВ��X"�7HY�&��Z��O�MZ��X����yF��YIo�׊0cdG�kL���Լ�LV,z�^�YKۮ����dc[�l�2��}���h��-�@!�d���C"�A�s����w�KǺ)�k���"�eK`�*F�
$��mg�I)�b��n*1(�������� uk��|��w(q�J;���A7m�r�W�_͘�a'� S<#%��?�E�$�%!�
w��)Q���yE��١u:(������ ���o�:�'N{�N��$m)���rhV���������r5���{�*��,��|�B0��n�=Y�v�~��#��G�������y�5�z�d��J�đ���n*���2�#��n9��k*ox��Y��(g~s�Y2����K��h���@�	�P��yKՒ��0u�\�e���\���ϻl�����L��X|l�����=�x�-�Cu3n ��ɻ� L�S%��~��I����z�����A@Nb[��s�b��8�N�Ҍ�W2�pj��`�j%��D,xݹQ���ԾO�H��$� [�jTA.��̬nCY(~�l���m?αbB6�w�rv�}'P*W�Da�Z�P���#� �e���(+媕�6&"p	�;B���䫫6G4a�6oaj���"��=����X��V[>��u�w:�kׂ�N���fW��(�HÑ;���@V¢�qYVq����g��۔�vo��ko����qA����篵��i�/Im�Kj�G�7�t ��T��C,�85��n�=�ύ0��w�evw.s� �(m�N�5�t�6��J�h*�(��S���)�����sB���B|ݑ�m�B�ۋTN�D��[gГ�ϐ��R�&�o&��~Et���j6l�A��ݒ���Ȫ�Բ�Ւ��$I�?s����i��W�q4�j&��H����}}\�&d�R�XH�@�ANs��w@�nq�wT�W���P&A��`%�{��F��{{���v�Ƴ�� 	{c���t/u���哔��F?R��=�z	���c~~�7�?N��Jt'�-]�tu3GNe��2%�)ብ
@x�ϳAF��=7����w�t�&�I�Z���r�{�|�Bi�l	��I��C/`1TZB/���N�-�����X�K�3d�8���A6ZL���Fo�0JG:r�i��k�V��w5����Hj�D����p�erA���6�rk6�e泫�5����[Y���Q$����&���/$�d���(âv��j�����#q蒚��m�}��;V?���A�����F�2�8�yɞ$PJ X�`(�'QϠ�ܡ�Ծav=uhi��=e��lC��Q@
��$G��k+ �i�*�/���v���r5��0gx%�LuA0�&���/9`����-[���Q���j�y�X/�rZ�}��r���5��;giޘhP�
@:�-�z�!�p�:��Y��)ӮV���N�tr�#��$�>u
����v��s�/���cH��{�F�r��Uz��2���,�\6\a����~*���8�#�*-��X���^~���^�g�f���&��k7�\�;d�ԷS�:���m�!@��Lc���J��Iҷ��τ�\�)�x�K�h�`{�b0�+��M���>�u�JI��>1�QɃa�����ؒ}(ps�4e�,�����%!�	�Z�����v��w�9g�^^��row,��R�HK�5�U�Q�9]��۶�o^�^�C���[��&⥧��[ƷW>�*cbjt#���V��cYL��L� �n����A$:7�N�OGh��I��T+�%�\>),ؠ����#JM�<ox�� �kЖJ�iL�{��~�7�m��ܛJ��f{n�ω<=G:Wf��q[��ed��q��'�-����Pn�ھ�)��G��e�#�W���?�R�j�uC�䀰b\k����g�"��Z�_�C,p�;����)�"��0pq[��g��j��[k���uQ���=,�Gd]�E1�/��3�����
بc�����9�L�ju��M��R��zԋV㾆0��amʄ� ��>1�H�1iX��u����2�W�W��v�s�Wo��%rk-<��N���FĊN{Kב5����m�]�}M�HGK�!^��4[���n�b��a���H�-�?v٦����ٞ������.�9�=�)�d�"l�����N�؟_�9R����C��]�����"tc��<��6W��سg�^���0�������:�R��e�׼�W2&$W9J�o��/�X{�� ������b�,j�2)`��ϻe���Z����)w"PwO{���.���`L5ȨK_4Ê��}Z��C� �P�=T ��Y�~W\b\H�"���/��Wq��/��!Y,A�&?e	@s����\\(SM�T`;������@k�/�K��j�F4)�V�~Q}l��+=�����h��@��B�I*b�7�B��$.3v�tv���p�Pʢ׍������jNa9�!2��9q��#*.:�	���X��s��:r�Էu��L[3���5���	F�6�D�c4o
I�r0�~�()�����X�.��7i��I�UJނ3� y���BÃ��Ϻ�#�rc��������9J�doz6Q&Q��q��̎O����`]v	s�l���L%vv��d|�g��Az�W��=Q��)<0�9A�c�1�2�LA��� �F	��H���)�nq��ˈ�|O�ޭ3]ę��qf�U�~xVqۏc�'NDZ�*:�l0�˜�5�J��y{�lE+���;y��r��z�ẵl�37��~�l�:s�;c
������I�m�Ѓv�
֐)�]�2bM��\�T�R)��U��bj5�o���i'M:Ѥ����s���2�	�juZT[בּ�5�1{���Q��k+�~����vVPխ_�zx���V3��,X��z��.�Ie�V�q%qj��ai�_��
�^��S�a�I�X֕t.�fQ��?˺���,�==q&~[��R����!qv����	1?g�͟&Τ5Y:l���~��M]���a(�xc݉�βaa�,�P�]�P>o?�L]���=)���}V�������԰�ף�[�*w3p��*M�[�c��EE {?�G!/w�rp��"9�ׄ+Dzb��F�e%���|���
�0 fX#��h~��uj�,6��=�����o����y5w���D���K��ƥ�u0��f����jÔ��~��� O@��K����+$>��|��}n��� wqJ)�}k}��p�����NO����}a��V���J�ڸ7b�+�Eyy9˩R,�#�����1MeF���W��H���+� ����~�Ј��[>KD Ӟƌ�Y;��rl�LKWs�^l�Hf~1�IA���%��C���g-��%ܞ�+�yIbaX���T�ЗO&��l�F#l:�C˝�	(�`�
	� y6�<ڦq�X������'ۆ��=�������QNF�1*W�]�� n�_��T�h_��L���u	��mI�Z�}�)��#�2һ7����Z��*;��qfm�_=�gZw����TAFݪ[�1{[�3d;��o!V����4��7��h���>
?�}��I�}�3����D�t��?V�.�lU��,�k^�� K����P*�n������l�_�O��$uH8�\�8�ߡyc���c��f �Ia��FK�37����&�j��7�`%���.Rz��(�㕃+�
#�8:�I�d܇UEKE���T���E�T�/��-	�IA�̤P������[�����{�>#(9�Ԕ�sTR���m�Qc{d�fek[�B�L��_���S��_v��h��6��������/�v��z,����\8��:�}Q*^UB�����*2de�$S�0�n��V�jr�$�1���G=��F���J���8V�k�d�L�F���7;�`�)�s�E5���[;�����:�'n@���G@�w#�p�!]�HyYg���CmU^�|x��:�FIut�'l�Lv��$Ӈ����+0�R�kO�'z# ~��ܜ�	R�H��ǋ�w�p�!���c�6��V`i��nڽg*G�]�vsl	�����L::�����fH�Xd�<�s�w��Oǽ���<��y�}j�[2 9*����,��E��!���!�G���=)Y������|[W-,j��:��g�z	>�a�E+w�E�I(�X���o/������t�l���Q�V��*���}[�\�"�sH|�Lr�s�~	*��h=y����~�V3�
-Ii�p���X��Py!ų�HJ��X	0������h~T�<(5��U������q���#>ayޔ�j�~��4������Е������X��ˢ�07r�i����⨗c��1����a�ρg��������P�w���d��fP�T�<���{�v=��ļM@��.0�&ግ���PP���[����L�aZ˙6���D�x��$���T�2�$��*����-Ź���A�1�Kr��7�h����6ik��:)�1k�=��l�S�Z�(��hEM�R�%����٢��K���6ە�JoPs~Q�`�	�;���I�P-��q��[��ϵ%���c.��$0�ZJǒ�3�ջm�\�~�Edn�Y���f�L�C�/�'߁�b�yK�!��X^\[6�%��@m$����k2(DR���u���D��K�*F�:}�"R��稢�l%,d��@�ߑ'/��C4�xQ�H+Q�u�g+��1��D,�F�1|
�n��qq&��P����y��VU�d�;7��e��(;�{���o��^���k�kT%"�!�@���c��6��E1��b�+;��m"#���v�$���㲄��
�j2Ы\�,(�������+�g����)z�i�<���Vpe�8�S�����5J��l�qK4��� �A%��;|>,jC�Sf�T\�/�U�*�Dҝ���.�F���aR�����U�O��{r����M�˻c��0�����Y��
J�@�Axvc��*t�f�RDi�����ff:[i�6����׷�ms�!��!>�@�ٙ�/'����{�P���y]��6{}��/`/� HUfݢ<�D|�cŉ�.v��-WS�*��ѡn���l��0�S.봇��|SqG�$f)���z�`�\J|{n�3pG�N�l/'"xW��4��}����\�Q��� �푺�3� �@���#�������������e�|2߾�G�[��0[t�+��¾������M��\���t�WNs�W��^bo��`놨���k�k�����z�W�����#ݬγ�`�А�p�tDTLc*�����J'/}�D&�����~P�i�\�m\#�w�=��ҫp�gS����C
��?���M�lB/�Ɗ~X�� ��Rѐ!�ڨ�p�>J�L�� X���W���xlٹ[�_M�1��.����!ѝ�N�����g�a������ �.�ڵ��T�[�Ŵ�AZ�[�(�{���E'�˽)���n�6���+cnU*t�JY/��ʠ�H6qP�RHe�n��{)ph�V�3c�$L��{�HA�!�9�us��G��O ��Љz�cLU�M$K=�ӎ����_��z��ѡ6�l9̞���}�%N�0_�I�'�&��8x�\ ��oI�n&������N�UL��}��%�^1A�N��)Z<��r�zb���Qn"aֽ����,�h�MQ	�����8�;)r�L�V�7x�N�)�l&��������B�|�v��$g��^�Ŗ՝CP�g,)o�fK6f��w�⠵�1~S�����(�e�9������`��H|�"��& ���$n��:���0|�!ɯ�+}؀�,��������-�^��������F��-����Z�x2�󊝥�-c���r�$��9�K8y`�p�\�`��p���:�CR&e�|�k�$�L�.:����[��:�����"xje�N=�FE��Ā�c��z4��mmf��{U]gq
�n/�ǆg�3�^p�'p��A�o�ߍ�\ �i��/� �)=o̧����Ƕ��u}����ʛ����xgj&c�%D�M�'�5'��>%t"0'V>Xcd=�%�JH9Dѹ[�� �\��a�;�A`Φ�d����p0yP�g���ŧ/iǹ̀��L��^h���j�'>�]A=U�:���迌c�'�j�jh�8�i_i�|������QT��0v�VD%�kE�\ȉk��̫�6����_e[l���u���9�Z�艫�67�^��!�G4V���d��e���O'��ƺ*2T�v��Q�
���$גۆz�̸}+�,d\���Ǯl���G��ƶ�+�s��Q�H'��5�rzA���nn�@󯊃�b^+X�mhqaCq=�T�������yRzN8��.X!��t���$�;�"���{ �?�R�o"4�f�3Y#�����3Cf�rm�z�)2US$�&�b%��\^�/O1(�v�˩�J��[B�����ж�_Q'�
d�X-��U^�Z��8������[�6az:Z����Pz���"-���	虢9����by��ȏ�#{:YЫ��K8��&3�6E@���9bS��,2���)�}��s�Ʌ~qt�Ȩ��#���_}��r����\"�\�FЕ�(s>
��T�RA��M�U�0�V7m^���b�"�.�����:��c�AQA��>���z�4��0�0_z�I��鋜�G��O̜K+�-=@�Q�X��.L*���:���M�ûr�qU��C<v��]�Y�@��ޥ�猀}�������^�(���b4q{�����B|��rl�P��� �#���ڦ��(hRm�v��R\�ūx��8�%<C�U�d�mV�����S¸�M���kSr4%���C����%��TJ[[��t���BD�{�٠�uWY�<+���]etM�孉3_��!l���+�ywE��l�2V/��0���0�p�[z�CW��C�t͉�_��l�z��.B���@�ot�)�J�����ɑ��-J��Q �lK4��U>Z��eu�[g�@6N��Z�ե)AOW��Jin�r���=t�jO+�e$�o����j�ÃGc`,�5VI�9��(�?\=�mE������t�Sa��
�	䵓���f��������gWi����u��G����d����6v��q�+�b�<��Xfs5x���C�_#�RI���D��Y�PSG�ۇj���Ez�I!�(�qJ ��wi�Zꂿ�Jn��"O��!�(�屍Ot���/6 gQ��\�=�#D���D���/x|6lZ��V��;"rؗ��G�V����t��?
������p�}��W���.��HK�AO��V��+}:b9#SW���#�`������vDQ��Pp��d�"����D��8�B2=Я��M������C3Ul6t�N��#�/2R-�;�u�&q�:	X�Kst���E�ޫW�W<B��DgU�X<�|�bp4@t�w�����Ş�F�gȷ"k7	AD�N���H�z�r�q��2�!!�c�7��S@�<��y:sq��Wn�p�4�ګ��k��,�9��7��1�h$C�����x�؟ -�d���/D�9 1O��:���;:�
��\ ����a�[(5��̱�����8���η��D�����_�� =(��=����Ϛ�x��$ �)����t�CQ�+�ߕ��!Q�^�y�X1��5Y�^�˯���d�	gwm�62�՛�jY�|#@\����3Z�Q2w���
����&|�N �}&�
���+�G���
��Pዉ�����2T��}�¹+��6�H������P{�<R4����������
J�S���\l�4 ��+^��<H���:��:��^Q��b�h2���61C,��A̚/��R��p*S�����t� �� C�	���3-iΎم����N�I�H{�Ь���6��SL����R�����qN���O�`K7�Ä������T��(��p��O��O-?)u������k��X$R� j�oM_���TX���'F&���n�@c�ܒ`��+=hՑe"zu��P����7.5Yxu&р
�O3:3����&�;��у]f���.M�[f�'d1���Ԅ�w>�)��k�@�O�}��?c0�rf �NkLBu���Wq3۪�J�$��x��2��õ��La�M��5O`8(*3�>���CxH�2��큶�4=z�e�i�0�)U�s����s�J��r�x/����R�x|ė��Z|�9f�������o���l>q�;�I}������������L���@��;�^}��q�_�!K�X,Y�u�3H��皴>
����ܔ���q��f��fen2�旖*���Qp�ŉ���U=l�~Ag�OYV���+��5��p�t.��w��3�� ����+�HH���4����{VC
���Jv�sA=-�ph��酙$,��e�"�%�)�]�+��;F� ��\��ԝ;Nȓ�ꊋ��L=5/Ӌ:�3"�S���g�����[ߵ���\��s�;��4G��ʢj��v�!��+����6ex4ե4��n1�bl	����B�%A*8����b"nwb��R��z�h{J��Y-mV\&�W�{jB;��hH)��|�ܪ�3gC1����y�L�k�+K`U�{����1Fg��q����e�����EQ�6�,(��ez��%�����N�:`��85�ﭲ ��.��QN|s�Z�w�
���gF۱���[4���\�2nU5�*�eyL/~���䛤�-��U�+��V1��TJ��tg�e�2	�B�-�˪�b	��^���$�'P�|��JT"O>��hb�ہ�����T�r��m"#��+ėy.+
�S��h�S�"s�s��M����Z�#<�0�x/���lO����⫏	_�O����ܠ���8�ŀOD��L�]G���#����U��M�Lx]���7�|v;qIwl8'>^r~�G �}�����t�dl�	w�k��a��o�2:�;�����}�B{�0kQ��=H�Bb�-MV0D�.����z���C��j_�퓅�jXQ���SP��.*QY���O9�׮Ӫ��E]��@EXњ1Z��]�;��2�1��) �ɭ���b�Y�{�yW%Pa������'	C�F>y�%����W�U49��D��7�Q�,+ ��N���J����] �W���?6l��UV*m�����c�W$G���:R�j���U��g t5NҦ��^�.��bF�F)��2"�s򟀭D3u�[�uV�e:�o�Z�V5�+�+l|���u3YQ=ք  ����-��ĭQ�"���$/���Ɵ�agE���<�o�-�z��@E)� ���]��N �e�X? ;:��d>]����_>I)R$c����׎t����2yj��fs������Ή��ۖߐ�J5��o8����K�K�%ZW����"W��&T���v�^��p���P�3U]p�_����2�xi�=�S��-c��D�ޝ`X���7�B�k���WG�V�C��Ջ���]��Gb+8�Pˡz�^=̻
��~!X� Z�����u)a������d�jb�����}�j�g+�\vF0�d�5�F%B�g6 �j�s%��R����V���
���l}����Z��� ^�ybV ��ڵ�Ѣ&����Ҿ!��/�33�*i��J���e0W%ˇK�]���q-��%�1���I���J�T�����P��Nz:[7&�;�@r#QU��;�ۀ����Z�����#5B���q��S�S��M%���|,P�Di]�KhJ_��W�y��\~	��r»���{AWЈlD�X���)���6�a�c$��`q^E�e�Y�����[ρ$D�/s<�^�z\�M�o:�+�][h�f�o�
�+��[�CӐa ����tQ?F�}���%���/`:�:[�:׫����o�7W��̞�7�1�R�)`WH�����a%�>{19,�EwH��o�l5��A���"u v(Of4���c�4|TIK�GX5�_3����:q<̐���2�d ��U;'z���y��A���	g%��H��<��:�4��U���;�j�G,0��?p���I՗TݻN�ԥ�u�AQM` �9�$"o��3J�ku+)1n'U'�������t��[��ٲ���6��2����4��u1x7x�&�ʥR���jn�0��Cf �OԼ�T^�^�6���a)G�q,�5�B�ڠ�����!Ga,S �"��r�N������J�'!�̈́����F���}�`��I|�W1ZГ�DD��kp��P��Q �ft��{t�bgL"�}M.���H/f�^D����#������"h�K�Xz���[�;N.��rƜI��;��a���CY����l@�� �z[�c��c�}G���J}ԡ��5�
B��}3�n�u9�R]�9pzCR#Wv��n�	�eb�MoP��@�`K\�Nc�.e`�~�`4�+��Q�=,x�fF c���5�i\@zY���%��ŋ�H����Q�m�i`.HY #�̡�6z��g��^��-��I�o�;��r��rm�o�f� ���e,���\P�F ޓ���ɣ��oLWΆ'Q���0�l��Rٺ�����͍7j(��뜤�C*��$�+��m�0��e��y��V�r�s�:$}��K#���ޙ��CLV�)����(�)O��"߄<<�߭h�MA��Ou85���n1��^��j�ףG&��P�E7�9�r����bf�/$�(4����5�0�;����;u�w?K}q5PQ�@Kg����,M�a��]'rH��w>/Э�n�`BZ�<��K۪�I]$�m�w�#cV�q<�O���%#a��g�m͇���|bb�r��U@�u���5퀃��W-���۬H�0C�-k����j��$C
�^�T�����@�a�ݿ���7�W��`]k�wG�C���������?a1�ha��Af��t�q9��8�L�QDZkSM��;&.*J��R.��@6�AZ-��2H�V�g������֍ �� ���UB�b�%�����4ؾX��߷k����5����L�P΀�;!5a4��jsj��E�%^mY4 n�\`h�RAY�E�{8>ʘ��V�j�+#��i� Ix�5��v�$�?-�F�/��je㱥�����V$aw����{qP�߀n�{a�C}����R�&N��;�6����0�?�hƬ�mN{oaV4����e�� a��UF?�zg���6�yz��KJ��촦To��+bL�������"���旐���n��U��W���Q�KL�~�ޭ0�Y^�J���߶)E�#��kr*SE�AS��ɗ�����[M�G�Ӱԉ0c(mg�M�ns��VL{��A6(�����6��K�V��s�t+��v������qQ2M�@��%2�0)zLS*|��� ˴: )ar�]���D���f��q����kb����z�}VJ��P1mNW ��gczDcYy�2�v{D�K�j��&�8WW}�{	ɷJ�@�*��?Ʒ���R|Y6�_�Ad\��x�U�F齨�yw��dn�!oE{�ղّg�--����}�f��F^�A�}�n��Κ3
@%
YW�jR�_6b���T��XcO�\T�I���=�%�g�ƾ�=�#]s��K���h�\��` +�[�[��6X����I!Z�Mq+���Nܿ��/k��JRN��x%��*fp�2��8���ۚ����7"�y�y�љ��w�b�Iv
�L
y����@�F�rED���G���O�~&�L$)��AC��m߃���=r���V脸�K�ӧ�qOfXGq��������?KԦC�~f�n���\��V���^�#L�*ؠSr��ގ�%4���cx
�<|�0 �7����m�p�
����}�ӠrR�~Ҿ��|�w��-f��N!�����qf=~�`��e D��gFab�r�{]����	@s?ۣХ��A@��h"����~��絮�2��M�!]��yY_6�/vu�>��L&F~�܆n�7��٘��7�C����XT��T#Te�{�r��_�-q�<;�my������]@��Y6��
P��%m�����P�'��i�Q"mWu��
O��s��9)i�
�����6���ص�eC�,�V����k�O�)wؕ7�� ~��"d�/'��?�`�9/C�ã7E�pE5���S5���}`���vI&�@>3�0�e�x駵��0(��Jk�nR.�� �qM����g�DN��"��x_;?��Z|����H�=i��j��	ŭi5_t*�<��
�Y���	wo8\��u�Ԣ<x�A6�]N
�������N�-�죿��Z&�f�{����*-�n)8���b{X�⋕��.�^��)��Aa]�{dP(����Ƌi�����ͭ��q ����}q�	eBj!�2���/<�n1���ʏ[��y��X�9����r�B��"�"�C?
(V�X���<����jLb�:j�����dh��B��\�݅'u��C��4h
���`��[�Ȃc� y�������5�5�<3�bؼ+�G����d��w tys�YZ!̙Ccu*!�qT��'�%�Z���J�5#Y�?��UiE�'T������!��B����BMİ�2�&0&&�{��*f��PZ�\T1S�o#�2%��	'�x7�N�P�!�~�3� ��Q�j��b$ ����'mh�n�x�ZY�f��'�g8�]L(�XJ�n9a���sq�A���$�;���T2�-)����0ކe��[�$�*q�xb��՜\9R�&8&6�ʻL�-,o����� W4f��:p�?�U��Yu R�7R3�r4iہ����5؃�k�a�����}�{�9�&��� K�"������;��{��&�}��c�p	-��j$�Q��4I�ć�
���ces��������ދ�F�#j]!$���V�qi���g���ѷ+N����TC����*k�t��A�W��:�'ʑmڧ��Fqlӟ�Kt�"�5���+s����
Z.PJ�cm�v�l����d�]��-M-s��}+�s�@��G��.���gD����h9q�ɥȄ�3�;�sJ&��[�D�Fp�{A�88F�#0�+}����q�b\ɨ�i]��]�z����s�<)0�Y�9ҕ��n�֛��	�y3%H�g��i�9�& 	v��V�����!����H�����󼦫A,F��&�����A~�}W�-�7Ҝm�D�W����0804~R��S2��k܀+@eL����2�9�n�e��M���P`/��\�����/� Z����6:Vl������_R�*�|=�_U����a����l�9h�-�`8�s�,����@�S�ಸ�|�"�]�OP���:����1�䟌`NΝ�$�)2K�n�3\.�>�l6'�j��Q_��yn��Қ5x�&�Z��lާ����PpX��)i
 !�%��$�|/��њũ���
Q[�mV4�99~[��V�z��6�pS9��h�����^��s3ꂨ�P��q[�4�e3�!_��C���6��P_5�4��#yQ�
.���C�	���y�Z���"0+���]�Mi��P�i����m��k�*�����F�7DIMjl	m�}�S�@�z�q�K��ȩ��Cx̰Tԭ�$�����#{^�f����6��L\3�#Q��4��Rf���O��#��:j2�����c�e�r��P�;B�{��z�����:�T���ZU��wmؒQP\pv�����a/᪃��6�)���]�6(���B��}����Ͱ蟤z^����jl6qc�Ҽ�4H�ɵ�11xf�S��f{�MN�I�Wy(�9y}>K��Ȍ�݌��2;�e�j��%�h�$W࿖J�`'p��������'FM�|!��5�f��W�Q�s	e}{N�2	���o������+]"1oϯA�2�3�#5YL䥸�^v��'u@��CK	�D�,`7��eE%h`i�OA�T�D�"c��.�J�VN������, ���E?��+@��4��E��m�����5ꃱ��ـ⬊}i6Q��5;�#R�bB.hY����<�X�;��:���K�9��~x�'����(�-E���<{3�4P�q8 ����Ö>�,38�N��]�������O3�g��kI�Ĥ?/Q՜̰��5��rǆ|T�;���H�LnW�o <�En�:k0m�Q��W&4{�a؎+hٓ�p��S�����Q��+����B$nsH��]�i݇oCl28��$�ʟ�����v,{�f�bB��&\�|�Mq����cŨ��A�H�tn�#p� �15i��n@�|P��5n���a]X��E`��Io�cWh|�P��)<קrz�B��&B�(.�l�,�Ѵ�P�Ҷ��	d���EF����R�bZ���5��Լ���'\���#�k�C�_�8�zWJ�A��=�'8蒮��i�Ɯ�i��_>��O���0X��w.L�;����0��I 7�$�sTS���#9�7��ؔ��b��r8��M�)=�y�T#FF�vG�/,BA�SgԈ��1�>v��)AP�nQ�c�ނ�˃?J�:H�����Ϝ���
��ك�\�L�7Հɒf�|��ŠX�
�����~�L��:*��}�/F�'	N7e�̽^��� �V^�<�e�>s''��s1���2O)I�y�}�%|`Wh�m�%dRF%���`�i�Bϥ�u�\H����.���e?�\߯#	�>a��C�(.��N.3�w�˗Mm���V,*�M�՜f%㤇)�c���3;WzOu�ڣ6��fA2oBw�-��a<f��s���,(	lM�ٍX�����j�K��@���%6������T45􁺓�ZM���4<� �G��d$��s[�1n�muL��#�U�_�kkJ(��pǃ������:*��{�ٔ���\�ފ6.�Hq�;�"�^�L-�vl�[&1G*^Pr��zX�3r����޺�C�U���ᴿ�����Y�Ta�M����E	4���Cx �
�]�W� ��}�K�g�J�����F��4'\#�c���'��c]�<�E�~�\bz4�Js{M+�gB�A�C�Z���7J�p�߷2,4'���V���ؓ$��W�כ�#�J(m�oVV����؜pL:�B�x�קBR/���M[(Tr�+Qp��,����g��(&�l0�c�=�d�R	^���ܝt���K�V�_�9k�
���)Ր�#0nB-	.����/�e�`N�急f-Mh�p����j'%�2L��}��{��MGLXF#���T�������t��x�49�����ToJ�)i�%S�����.� �g/�R8�s�V�>9�
�ߓ������]�%��9�ҁ�����ֱ�I��� &E�4F�9p�c�x�V��(���)���lg�]��!lQ�q�+#_�a۰hD�"������:�WgQh�ܞV��FR��0�d���r����)��O3m��8o��} ���jW��j6�9�.�\j�ӗѰ־�cC�s�p�	��9���m�<���f�9�~��j��E��&����ca��ź��� Ճ&�^h_!֪Y����􈈜hi�������Í��_`�&S��|rĄ��r\�{3�C�C/��acq=��|�a")��pA��J��$�b�%(B�B��<���?�j�ߥ�f;}-�63��c_ �B�6����śr v3Q�%z�c�`��&C����źa=�a��̡���(��M#RP!�2T��"��u��ԛh�째�,��,wy|.�,���(�H��U ���~s:@H>l���[����nK�q^c�v��x�l��N���` 7LS<o��J��K{����~�'ɲt>�Y�i�X�}����~��U�=�ˀf���-��B�]�k�$y����(�D��w���:�`����$Im6+�̤�'~u��V����?l1 �]�h҄칾��s]���#����\*����sѿ�j@��,��@ǸT�<��EI��ѡ�?!V�9���rJ.�(8{�����2�J�"=��rK�����^&�F���I�G4�?�Z���0
=�"q��y�(SmBQΩ��7�u^DN�G�z-��s���^����K�
��R����s�P�΀�֚����ty��训��S=̞���V�^��s�@n���VD_e��ɽx ���>�X�}�=��J��񥟔�'�S����Iqr6v��9��_��=3���;��fa���S�Տ�-`HOV�pJ΅��|��W�C�B_z]��������/zYR]g�uz�|����9�-�z~�#��B�=�l1ի8�a����N���d���)�.������!�F��cu:3Q�"Q��)Ka�\�W�ȩI���5)�!W��2K�:����55��f8d;����J�O�l�+eUy ȟa&.��,��.�yvSL�\�?B�����֑|R\v�}��G�t�
�<� ?�ņ�^�(6���f�]b�H�s���W����]P)����\����*;�~�w�3�N{B?@��9�{�c|#�:wQ�����@$xy[��;,��K�@�����ê9N)u���Z7��h/������)������P;��L�+�����Z���{����i]�0P}ʥ�v�"��~�6F�x�£,t�i�st��Լ\��m�{�F8���vucҾ�>�K�f26E�n.�[9f�p�	��m�8�@C�﹟;��ŕ�ɋ 3�j=�����@S��eGG,�5B�T���o�ł��E�����2���XG�IaD+�Ӭ�
�U͙��&��Z�`U��!d��k��ODr��M���z�M[&���\��nO�htf���<ƀs���psr�i�3��?3�dwEd��0�+,�}^7Ȇ�\�Sk����=Vi�qv��z^4��o����~�Ͱ����s��s�)Rlj���I3֦>�Kz�WE����gה5Q<bZ8
��Jg�ְU10��Uߗ�C6�p��9����F>�%fVV�p�0]�$����k�}���D�
o�I=�ɆYb�y��50�gc΁b�3�z�ɤ���fF���>�Kaaz���"��Xmo�6,����Wi�~�D �5'�H���FA%rE}�������P����3����g��%��f���lh�e��}.Fl�4`�����m>�AE|�l�{SО,e�ţ�\�����Ͳ9�p�!�5�(���^k�D���r]|..3\�sn�d_�E�7�%�*��-?��Uq��.2l n����f�[l& #]�]f��S�W��	��"�A��P���Xgo�C I70ڃLu�|=�~�������"�t|铎o�)��wO��ı���k�~��]��x8���T{�p�hO~Wآ��M��)կĩ7��b���se�a}�[6�>��(k-d��f�Ru]��r!��Fࠋ�u�q�z��� 2�e+Q�!<��ͺ���S�{[��8 ��ĥ��}���.7��"�.�k+5�Ξf�������$-.s���F�ȧ4i)��ʏ�InQ@LA�2����UcK|*��2�&{0E|����;��<cRv	"xlK�ǰZ^�>�Ɉ���7ꕚ�#h�+#�}�O����+��pF��^�uy�P?�u��Ϩ�w�1��ǜrS�	�,] �:D��$�!f�xF���E]V\���s��h6B���e�A1
�pʵ%��.凋��1��`׵����|$��v<,`�8��!�;:B������wܻ���S��rT���|o�U&Bʹ�����ϸ�"�N�ds$sX="E2q��8X��_QXi�%g��=��Z<�@��Ռ�g�f��K��}��Azҧ�(Lv�ˤ�!��9���	���KOO����I�)�y &��	L��;���NP�"����.�^���֒��	���Xtc��N�X�:ߕ��sIj�hy�fs���ہßl�"]��$R�I�;gB?zU� 6$��B�T2d��9asʔ[�;�(!��b��a-?��9�K}�yl���38[q�"�|0������/N_�q*T}~�Z�FT�r��ʁ�yx�������:��qvs���I���ͫ��e�Я×�^�62�I4D����V��e��+���[�zJi�(�e��r�m�澘�J!
�K�?�2
�+��%�q�ro8���Mu~f�ln�p>��=u�+/���CRP�J`?B[mja�>��Z��!� y������
{:���8�ݣ}�81	?or2���5iM��ε	ؠ��^W���59 VpU�G]Q��-b~�0m}ˍ�*���Z�~F�,u�IG�C�hM���F[E��vD;`r���\?��	g#���9� �s% t[��sLjl��Z�r����ա�S���VF�x�1���Q�Þ��3��Hx��}�d0\�H�Aq�`��@�N����!�,^�وՀ�8#54h� yya������p9�*��9k��-ON��庠�4��* �,������~1i�?${�e]�Ux��6��:��Nl�	���7ֈ����xH�s_�"/�k���5���v˭YU{�yD|��&2�R�7��>r8l}��{����a�GD������ ���7qmY�ąU܄������{�V~�(�k����g��ۂ�1����y���ЀU����G6?!�S�^�@���'����W���������]�a��V@�ڂ0|������s���ӄ�3͗���Tf���,�#���֒=�Av��"��k�u��'Bt'���CG�Ġʉv4��4�%]�ҵd�ib��!�����VE'���*Bo�cR�Qs�`�����"��<�E��(\����B��!g �Б�s�v;UaԘ����!X�$5ySxaF��f*����#eMݹ��,
$\T7-�)��u�V�<K��#ĘT@u�r��	:���[���NK����*/|�G�UN�s(��Ƥ��'�LUL��:�@��E:ι�9R�^*�"q@5�����e�H���G���;��/�SWk(R7��(>2yk�7��.�^:�n�EՎ������o#�4�V����0�ۘ��%e�Vu1,��?�'���t�?���l�(��'��r��Q�?��^=�8��j~���x�4�^��
`��x�M_~�ڂ2X�Y�.�M��`�@�Yk���}h9��0��"1�,�d#vW|���1����7��R���������g�3�w��(�I�`��*��d�˙�����F���#�Py��e���r�>���A��}j�,k�0:�@�>ٖ�@m
�o!������[��e�j���р�Nz��-�U�n�ފD��w�J�w|�M����J��vr˃��C�T��A��N����] ��R�cv��)����Ç��C�
��摢�:~I�a���pV�=V-��'-��\(�R���r�h�b����#����`���=��ujp�ǅu� (�0�����Q[�pJ!80��;ÓCx�X><��E.�r7�;u���c�X���G�yQQ��-��R�l-Mn�|�?�����3��*o��'mG�as�}�>���L3#m���p.kz��G����z1Z��wS�I�g���|�0��U �TNlP��x�Ih6[�Rbj���KI������I�ǐ��0k�M
�-a�Nt�Ǔ���kv�9B��k��Ni�y%�3��ё�S+�w�������uCÏ�ٕ"�!+X���V[7�G�$J��GX�>�bo�!�!`è�MF_-�#�
L�CMJ.����l��g�7O��1kѨ}&���i7�D����K��f�f~*��^:�ڑ�M������ς��@���	�>o�����	�K�=I~ʀ��j�Ld-�kLHd۱��/���Ms��"0]�Z�C\�U��1˰�d���q6^�P5 f���T@���aMi�n=��
�����?n��n��5��~Ssv+p1|��v��:@�L-���6:�/�WWF�	%�z�sP��	������.2]�N�	��͝�j�6X��=�=�ut�ef���C�oeJU���5���h���Y%�ᘑ�gM�&3���%�$Y�����6��T��- 2ȍwݺ@]A�S�%h>e�"\�c��Nfe�ͫg��H@�h�� ��'�>w�rd��Ԝj��s�+����(�`|N��|�sh��b1��ֲxq#`J[O%T��dRU1��q��(�)!R]�F�#�2V�%�!�W`��7Y��F��akϏ���X5��<SǢH�v���nmNx���6�m>]�e4���,LƢQw�6�4`yT\�o�WO�.�$��"���j�b�Jv�DAͿ[�N߇�w
�����Rf|�qalb5��6�y}ճ���^�ذ+T�l�9�a$UҾS�(b0�^���ɏt��㧁�VH�篗s�~��k//���}T.W(g�B���b���H�v�8B{�i�8V`��'
=��L��G��O��ܩ���d�m��C�ޖ�@���2��T�F_�ۉ��{��Y�H'� �x?��ns-��)��	�&���D�O>�k�]R�;K��.T�d�R��.��}Ho��cw�0 ��=�w���QM��~}�!t8]�f�������1<J>qSD�і��`����q��9��R1G��o�7ُF��wS��8��t���}�z{�7Gep��[O�9��zm��l��� Q0v�XH%,�"���K,�{�E�aS����Fb�y�l�(���q��">I=_ e}d������o���������~�
�	1@�^�N&�<�~L�D��f�*3�z�$u'P��A\A��q���|���xE`��V��i�e�.h�<K/E�YU��
�C�;Fw?4 ��6�i���_�gO�4��:���0||J��Mo�@Sِ���7�#m�lҨ�nfY�} �����o��~*�o��ăਡ��B�x�K����=�U���"b�|m'rϹ�si��O���G7'�	�们[�R#O�h��f��it�ύrq���y�
�c���8 ��@ش��n��5��ѨyP����|J�S��� ���;oȜY�S�淬UK52��	���@N�~i���b�#�隗FCOF�b���@e&t�|���Y?�X�����X�,��_����?����������R��vD�n�S���ݑ�7t��caz�+�ש�=٤/���{�#�WF��������1.�sR��r���}�x'9��� `p�#��f��O"�~�����jW��{㨺ϐ�	��m�o��1�벤q��z�e?Ւ�Я�iX$7���&��������}b�,��wp�89��q��v���J�:D�jF�U@~��9xd�\96|&�}��l�!����̃[$��E}a��ˤ^����^CfKkH �=�+�r嶻{���[�������Q��V��
��N���Ͽ��q����xh�H��K���NN�+��e��A�����z��EV�Շ�|VCֻ�#\�$�?��0#Ϩ��m'�fC�B5[����MaU��`Y|��M�P,��lՉ[�Y����}�"+ik����9�-[<�V?�r�d�E~�=z�P���2��W;�N46�H�Y�Y�W'@�9?���	n�I��2�Qw-јʭpJ�Cc��U;J���!�ȚW?��q����Ye�6݄��H��^��'��ו�7*qm�@���5��	�䋠o�t&�
�NРZ(!>6Hx�³$5��ɫ߭`�譡��Qhy�R�8Ũ��^����U+ïj$)D��Dn-3�jt��;��qP%X���ع�<ɱ��KoË�NP.�7�$(��	������1HPw�Fl�Qq��j&���'�4������/6��W6�(��+Yq�����?K
�>��4�;K�a;dyô��?���1�����rJ4H�u��xX�˾�ь��K����h�~�m�0��R.ZG�Ϛ�ۈY�B�T���� w��zpZ�\�-v��|�S�&k����\;�	5�蛠pH��)-`��M�e��&�����-Q%��˅�s(��}��/i28�tUk�ԭ��n����d״��#Gd��O�QE�N��.������o���Vq��~�����@�-��j��>rN�G�K�}���۪�
�r~A�&@���VQO�C#s�{���m�t�r��&�!���W��Jy�Q�%Bț{�={H}G�W�u��e0�H�f�OeK�P�ͿC<���o0�w��ϰ�m�5Q �=�J��(4��ډd����*�^B�;�G�)�닍k�ӘX�c/�T#��K�3�KU����0`�?�=�H�2��@?7s����K�n�\��� 4�˳�E��_5^�/p
֛H����T��L_7����n�6�׉�l���}N�,s�$�-՚�g͵;��}9���\��x`r���i��uw�c`�V�#� ���̊�*3�]��ה�R�+���X��h�w��]�o�P�D�6�����o G���g_�6C~�=�Z��&��nT��q��I�iꂄy���ZZ�.K$cDj:��ɳd%Վ��P���:+�P�2�j>���9�E��-/Ƿ|�I� ��&��~�x��c+&.*��s��a�^':��x�X#�3�^��9W�`?9C�,��c�Z'/��*�c��9yh��6D��6߂ʺ��No��T�	��n�8��;܂Cp"���Db��[��K�Q�0pqS2R�x�e_���Rz�d굦�{��cr��@ �C�r~���Ӱu�Y�A2�ة-,z�	+׼�9%���h��;�;��|����پ��`��O�@D��M���|����ѿ�RJ�"&=�����{f��I��4I��,Fʙ�#d0r��R.*��>����7>K�xz�_����0�`��7P�H�m�Uf�^��R���7"D��t�A�@�9~�#�^���T�Ur{��O0;)�_9j�h>�P>�
���C�K�{�x�#��svd�(�ԧq��W��3�.L�h�{�[,�i�="��YS����N6�~�����q�H�2����[��[�!M��e}�E�����=Pw�󐻄F����zR�g�f+��{�Xj����
�-�>��㵗Vrқ����"wn��#��F�aK��!8@~�9t�>�Fk��mR������w���x(iրX����(�AC��9K�u��:ַ|�s�m,d�x^����0�[�[iQG�
�o����-󢮎{�x�F}U�ri5�^S��,QUXk��X^�q5�������
�`w;�e��ST)n5���s�f��h@���$Y|C�|q�k����:�>OW��9�-/J�r��
!��c��:,fʮQnt���k���7}�9�(�b��4�׾���f��pdU*���7�'$nN1��Yl1�r�Q�������(�U?��/{��X�t��T�-��m�F�u/)ㄫm�=��fX3��q���rϚ7(q�D�.LV�]���2υE�pb���8��c�ruOzѾ=S��n�}�	�V�=�l�������,t��������<��N��	J	�#�����2@�G	[��*gu�P^IH�P�X=�^b��
w��B�������
Kve �{�JXĴ���v��Ho��S���7�缔\\h���������e��O��JWmt�� ��'	�I��_W"��O5�Q��	ld���6@7Xz�0��̍�Wf�����g�=�)W/t|����*f?��7���t���LE��?��ʱWZ��#}	zqUݟ�-3N��+�3|GːP�[�X�Tb݋i��{�vG���jp�G���)� eR��.���i�`qt�5�bꡣv���^�c�A��JЉo���O����6�6c���ѿ&8#4�_��� d*�sA��1~�$�
|[L��RG�; q6]�$��3	T�C_f�ji���؄�у�|����Ms��J�R�s <���mP3{����g^Q��p����p��We��Q :��V�0�ߴG��c����$��^W��zσW�Ǐ��:������յ��1��,����kS��{�2���A��ħ:�w<�/�~���X����ӟ�W�^O�=�R(K���n�c��U]���� 0�r��<���U��7f)R��3�>��?L�}S������˃Ɔ�s�q�"
���P ̲�]�m+��!�=���=,�8%�(@�F������S0I�5��[��5�A6H�����DfX����$ϼ�u��4��2���T<�%�$�[�˨� rW�����g/k��|�D��6w�њ= g����exAH�!�sB<���o���On�m=&Sz�xaM�ۊbj�K�dڇ�|�q���|��1~(���}TF̀�n��e;� ���M��ǜ�!�PR%��Zn-�J��j�� ��������Կ�aP<�� ��PA�]Q�jja+ѻ� dG�[�����JE�5�1[7�aD�ֺ�,��֊b�?�m�y3����3�o��T���$�Au��.�pt��q�9�-Vʿ^I�<�����t�ua�;�����6@i��BY��xq���e`T¨���v�O'�Ѭ�q�>o�P9/96���եpuDU�l�Fi��)�oE*j�lf���e~�[Tv��$�Q)+�k�)�^���|_��_(E#��AR��堖�C��/�M�n����*���A�J��h�.����w<���=��8Q�t����6�uQ��rS��J|���Of�k=�:�})</a0fߊ+�
|J�h�2B����&����囲vyL �v���k� %����������ݍ��Oҗ-ɞ@"������ӳ�����"�<7��kf�sgVg�I$�b��(����"U�F/��V�	q���<����q]!*�<�8�8���Fs�j�].Y���ry+P1$/>{Z8OJ�mA]�(d�(�����������Z.n���L3��r)@,( ��0|�����r\��Mħ�γ�㘓��~CJȺ)٧��Y4����s�¶ɞ�������}Շ�}�~�4ac�=�V�:?�B9N�}����=��C�&j+���7T���}�����'�6-��Z`�C0�Eّ((�����WD�	�c���$]��7��&��i嶈�u(T}bP��=����{[�&�U;������uqo�{�4y� 9�xr�P
��pSL�ڟZNY��0J�;[��A����m�|竺�q��[sU3��,�����Dox�F��g?`L3�#|Ni�����.�+>�M  �p�D��C�N�]3��!�?��l��c�̮��_,~��u>��ay�����G�V	*=g�N+��%�+�P��>vH .�.n�$D���E���3q�pD��U�L{r�5��֚�cd}V�u�ʠ�����|���!pSk͛���b��A�(W�3�z�w ΃��1��Hgs�,?�YIw���Rb����鵀�P�&�S<�l�	��y��D_u��M��N����f�w��k�Kvu$���Ȭ���Q��ǎ��yy��hiA���H�jՠ�����7~�qz�n�ҋ?}�/��K
�1-$Nߒ82�)Y�8��|##����́zw�l ҷ��8g�cs�#,�����=�����}+\�4����Jwm���?1NVO��C����q���,�ݺ��0@�����Bb-7�̔�N�7˾���6s	�ledË�z@`=�'�_�Z�����[��M!)i�m�5�{���F(��6��k-HX�2+���:dN|CQ���`8�j
X��Ƃ�����g����0�ш��U7Y�]�-�Dځ,����q �>���B��0g�i�{���\�Y�S}.%����q:h�'��w�-�~�6�?�7�g�� K"���b�b@��w2r�.���5I��o�y�ÕnE&!���[��kZ��~�N>�h�5�Υe��e�7B v%��J�>:H��`�s� $������G���E>�̓ĵ|���f��R���p�}$�7&�Πqł�t�C�4�H��4����+�wO�c����h�?���V�5�g&~��?U��3��s��Ǒ}�)J7�%�wY�U#?�o���`pXS�fhUKk�-��ތ��M{��v�6:�1L�*���F/�I hy��+z�HJ��o �0�NV���Ɔ1�E����]��"����X�i���	\�ze�����;���d��j��H�d����f�D�.�� �]qM����������-�S�$F�B���}hK*�6�yyd����)�<ɰ���nh�(��'f�P�ܙXk�T�߆<8��u��Zx��l=���H�Z��."/|g'��P{�;�HDփ�� q�zkjtק2X���ڼ>A%�8�zj)�P��E
c#.x�W䄞C����z,m�/�>P���^Qi�S�^��|M�s�ݚ�3v���&�_g�-�Hӵ�0d-�zӥGa�U�/I�aLD�O�k���� <�X��8�po��E�$u�hv��.k�i�|��-�9�#p#t�q$j<lsP�q�*>=��mK��@j�/5�)*��ڒ�(� �7�R��k�:�D׿�����ʎ�j���}]pδ�Y�uY�gO��j���ղE���]QЇ����֩��K2C6��]������LGSQ>�Τr��S��^�9�d���(�i��9�M7Ј�$\����� ��<��q�U��t��Ҽt�9	0�����w�9eH��A���@�$ۮ#�I,�?��#hq�tHN{#��WP�6;K��-,$x���ű+�(��JDЕ���� ;In�F�mA8K�,r�@���B���e��f<�*�X�m�N��@���M����4��C
���|%�ٚQyN)�ݳN�i��O�ѿ$�-�5,�T����r��Gf��[�x�+����Q�i�2���:�7DO^��M@�`d]��T1^����96���_��5��(��������?�,���C���@�E�Ē[
���7���e~�T{	�%�JE�W�,��7�j�͋�-�sO3dZHS?4�	<A&<e�̪��Y����Dph���K�ȣ�:���	�aw��A�EQ:�ؚ�4�jfQ�K����מ�� ����_�\������9��^a·�S��R
�/f\Np&G��|]�6d�D`g��:ר�`��*\{]dܤ�Y;�� �C�t��`�����P�R�%��M�:dL����{��pd0�s'��g^�	5_LI3��s�K$�G�܂���;#�yG��_�Kٞ�捎�Cp�:�V�#x�:.��G�,�1)��x��J�j=��I4��\�ޭ:`�O��BZЪ7��c�+`u��R�񯑶<�)2����?�!I�
)���^#��w�us�.���
L��\h���8�Qȫ]6�,+U0*|I���ޗj�f�|t��r�CbΌ��t~#�+�n�8�.�r48�n�2���²�\X<��`�A��/a��y�������pS�p:� �9ZNS\��N���+��P���<gV�/LZz 
��p�v�AQ>�]�؜η��Ĉ)O B��hx���j�>\���a��\�'�i��݁]#R''1�3�X'����#5�LOW��C쓤5�|�'���8�.#F�b�!��?êQc^��~J�W%�a�ٖ�@�s�P �"�HvT�"���f��%�NXs���. ��Y�jiJ�j쒴�C_ 6��,�~�s��e3г���ź����4jl�\[�0B��R� I�L�BņP�6 "����+(<Ĺ�l�<�Ǆ��
�����^�6tUS��J	����T
Z���g1ء9"�^RS�^��w�D�&�����K�,��]q��@S*��A˸��k{�Ow���ԃ�v��x�4$�j�R����>���������m�:�!��T�`�z�V�B1�AL|�^��~#���m���S�W2�M��7�3�	֡��3 ��?i�B�P��j,�n���Qg��2I6Ț�E4��W�F\���q�@���l�F��0�ӎs��[�C�7��G(����IĬ�b�;�G��-�U�C���}��C�
Y\�$Z@�;uOW��٘�Q�?�	�6EK� _��<4.u��;FhX�?�o��gS�Tic����ru�)�j�7�,[��ⱑ������� ��B�Q�'��^�G�����BU�� �l���>>4�J�s�C��cE�����(�
/���{M�θ�Ѐm)�T!�Z��l~�>'ٰ�º�r����.��'���|%[�J�p�(�#��'dU3R�g-��,9X-N�d��wQÄk�X��3P���ۍYQ��q
P6H���u_Pt���FvZ,�?6���<)՞�%�|�JG��G����Q�#L�x�c$́�F�BR?�vFX���Z��sG���܈����n)4Z��������h�c�_j����1��7r�^oGڠ+�)���xt�,!���Wc�(4\��G��t�9���t�RSnoeL&	x$�*2�����
�}��+�9�^�%b�b�_1(�cS[�n=�B�n� eD������[�U�.��=x�!fk]�[��P ���yi�F�#߄$,�F������ΗN{2�����>8�%�=��c�r߃���v!����5��q�|+3^�3ZV�-��X;M�+�
��Ø�w1�"02E ߹��T�����e!���Ԣ�٘�o?�o��u��yp�}��σ�ֆ���R�O��U��s��#�4ԀG&{�}��%/���+A����k4��|����@��6d�Yҟny<�� ��$���������+R��7�1���(�|�T�����G�"��F�ef���Q|v%�'�;7p�|��f��k�c��9RW�u��Vh�?Do�%NY����%��e��oc[/@lBy��iy�B�MІZ��S8ӱA�e��7�����Tn�ڹ���.h�,'�!;C�0<;Q�y�(���dz��,V����J�>g[�P��];��=&QSn�Iϼ#�.�S��c���Sx��q-�vXJ�;�* f��P%%A$a�D��5u1�1ʂ�Ms������������?|�C@Xm���Μj���h���7]���(���o@xp�I9�71�|A"1��7"�p����-^�w��7�Ŝy|_�8�tfqLw���[ќ�9u���f���u��ř$�E�i �����Ē����8q�2����/�,`���8I�,;::����ѥ$+�'t�*߮�Y��P�[;�(�cT�\��'����d���M��I�G�+�d C�#Ԑ%2��O��_8��é��j�Y(��_���+'_�����
f��u�N:Uë����Z_~}� ��Sž��䳑yG��C�e[�־Qn[�_-ҁ�Lh4����d�05�*���@b�Jϖ[��{a�@�>L)ܽ�[����`39E{���hͥe�������0x~��yl���"3���p40l���	�XKw�G�ډ��=$�{��ˣ��]a��M�0�_K� w%�1�ct��6����G<]v<����ʷ�␽�����w1�a�Wy@Q��w��=�*� V�]QA��g��[�n��A- A�K`2�j��3?��f�	ܻ�;c��[rb&1Aۈ����?��R��t�?�20CP0�D�^��c~���$��Y52n��g>/.���!YS��F�������QzV���B��YU;k���B���a{�v�����Г_�n�`#�䨫��}�z�E�btlevm.*v���l��aq8tJ�qJIO�txgN�h��9+v�������﾿�ʑӥkM�i-�sg?g[>�Խ�q�Oc��"+n����l�< Q��L	FV'�o��J��%�
Ƒ����!�<k5<��xp=w�x�)-F�7�I����O�&��򬹩.���U��{�U=�߼�˫�r�ye�Up�3��V����fj��	pL,e�q��F<4�	[7���҆����"����mYV
L���P�.���������S�)Կ�:�g��i�c�s�<�lE��݂��~���M�����P��й�	�*� �%ް�ƞp�Ŕ���I���Xn�pV��6�N����#��Gn��K�6~M=���:��E�3&�e���pQ�W;�-(�RHVY�xn�d"DNU�x��W2_.4�Q��K��T;�ߡ����Zo�V��DˊG���z�nl�_q�daZ=��-���S�� X���*fOxײf��٭�I���O��9���8%���ku3�H��]�Mc�5�<,8��D�K,��%=�m�~f�+�x��R~��"s=� �X"�98�KB* �����U�L�M#����@�
�QW8+��Z����Z���vy_������d���gc�N��2��!�x���4���=#^�}���ˋ��S�P�HgS��v�^
�[��+�đ�
��㬄	�P���nm�4!�������
��4�H������om�;�K(�Q��{ o�ȳ��ze%��F	��Ȁ �|�o(����ϴ��Y����y�k�>���1r�k�+��� )����'���6 xxr(���n�G������Ȃ�%57��G�P��,;����U5��q~��g�k0QG��sP�WV~����o��)�tQ(t7�W�/+ ���e&�y�e�6����I��pW��U��m-��
�V�*�eX���MsE�aa����Ǿ�o'1�x�Z�z=5BO�z l7�g��d���u���M.�[ IǞ'�Й��5�g��m��VL�&��CRQ�D!�R�J
�ݥ,-iƭ�4@PN�8�� �c�@��}o&�o����Kܹ�F~b����];v���g�5��a|fQj7_�p�\��7�~�����"?~�u����.���?��(���w�!)����xP�$M��T�u�-9���$f)�[��O�k;������-A�JT�`:iz��UK��߆N�!�EL0V�C&I�s��ODoD��&X�$��e��l�)�c�_aC��3��ߌ17Y��2U�C9Tj�B��G�/nڻ'cvB�X�2�Q�R�ܗw��@6`g�#]G,#2Ğ�K�Z����MR��v_l񥩄> fy����K��5�E����5@��"�޶#,9�f�\�1=+��_�d������':Z�I~�|Q�zY�GJ�z)���^�ٸ���vՋ������[�e�d��m��"��� ae5��h�:��Q����o^$?��0/��on��'���Uņ���|۝��5<l{zɷ������C�l��2_e������`��r���%�%��}]7�#��QQS���2O��x8��A���j-��-�Rݑ$��[�D��2��\
;����+A%l�!�|�6,���ã���硓��[s�J�@����(�eY>%g����*�k�0`���L�3����}��5�1E���ӆ�k3��:Ǒ���緼i����Rǿ��� �#ae�A��$_pB¸q�£)�S\�(m�M����A1�K���l�"n��v��"��4���u�����<�m�
je����)�Ꮴ��cE �R��芬��d?��������S�������\���22��˔
�fO�9n��~z��>s��u/�YF�c�P���-~��Y)
w`y^5r�6�a�}��{qv%��]"u�]E"���
������y3Ѐ��J3콼�{�� �H��5P�O�r��p����I�\7L���7�,�����y��H�]T�p#,�]��Qn�mUV�G-zq[�E�kb�b�jBZ��QB�0��Y�d.U�L�=n���i SՎ��5y&����E|Й��=��y��K[}��yh���fK���g`	%���)d�>OQ�?�h�C�wU�A'�C�� �>�XkLc�uZ�����8�������Ȏ���]'�G� 3�����240�KQJ�CV!*�e��g�QrL�2*\�k)�zT1���2Au���qK�1��\Y^P��T�ׯ_ڔm��"��|��%dLeU+L?Mӱ"lb��0���+Ds�����Oo�C��SY8��WPf%�%�qmӌ�~�k��Y��
P�M��Z>��2��b$<$��W��#{�6A��Xa�l�S΀D<MYUac��UU]��Pe��@�I2�>�]�se{�T!E��l�`��f�;v���c�����@+Vbg�Q(���nn-$ǫ��g	����*�miw�y�b��(���f�R�����w>�C�ɫ�~Աӯ�l�u���]��K�F��<��hh����n0'_�3N��>���b�?R7��$Pk�VB��)���~,���lY�A��w{�U	�{M��+q�룥�4B���Ƣ�A|�����u�b�̧%���:2T�I7|�"-�>�1�C����]<ȯmG�(\�x��F�"�bءW�=��S��U7�1��|r4Ii��9���G��Y?,�]�N`�����oo"Y�������Vj4�S�_m��i���h��K���=��~��tq���=F�=UGdu����	�$ת�J�hv��i&r����,����<���v/;(�-�g�h��&��O��"w�o-�p�>��m�1#$R����4k3qx��=�yUq�P�<#�����GD�Z:I��a��%�q���;�I��q]�1:F�����$~+z��Z��v]����'��&3�f�
�`�{�9{,�X�ʑr�d]eO/��D�P�+b���q7��N�T�^O'�۵��*o�A���nτ�<Cq�����8c��j|j-	��#��R?���]6�zj�L1�%�j����w忱�
6�GY/�	�I�
���<�n�i�
Ib=C��2,p��3�3��=�q�[��5ʘ���p�&R�[�4��l��M�u�T8]�c�`);���c��$���X^9f	� iVx���6Dl ��D� ����[�m��8�ވ�7')z���q�!l�7h���,���4O$�z!���]\��`�uY,�g/�/<��";���B��1N���M��s%�u��w���J��X�M�z�,5�xs��@����I���`ds`����6�>?�gpNω�L�kU7�x�_!�buO�B��u'a
<�+m+]#�q��Gk����:��|��?ċ��6�.x=5r�i���Z�����n���(f΃����O��W7��)𡊲wK=G�p�X���P��yOTH�<~���sf&��i�j�ct�|�p,�4����,���"$�t#�^���N>L�=�+ƜX��?w�"�����i�m�SEºk�|�FDC �hK���`׎Yż7o�^�<3�I>�����.��+��p�'���Ѕ��Ģ�hG@���,�9m�oh8*�^�� ��	���0C;�Ǭ�3F�T}}�i��.�Y����.��{K4=���`�x��*�����D�k�V�!(��+3��#���k��j�I�H?+�l0�Z^�~�j\\c��.�`���U�W�C���k�:�p4w��;�H��ƳX���iZ:dÁ�h��c �BKj��Q/��ՉA���:&���.�s��v��%����ٔ�Y߸��UGɡ�H$���)�k���l_�z ᾯ�Q�c���z��%^�$ �瓄%͊�8X�r���L��_Ed���vX�일w���B5�.I5������ D��}0��v�+�\�W�-:NdF�]e��dh�Y����ö�b��gk�p�+�q�q��r���%Ar! t��'�n��p��D�Z7�:0�U���wB.�V�(��|ߚ��J�4��y�2���7��`J���U�7��.�.�%_�;�#�7�ʑ6JFe�
7��O��h��VY\Hx�f# `�u�n1n��K�l�w����_�'
J�b9�U�Sת����N�@^���E�1lU|`����� ˠ��Vu��d�H��h/k���Q�1��b<�ί��V�A����j���(@g;n�r����B��V��TNsm7��21���p>����e�?�T�� ��K�I�9�����f��S��,}�GS��^PkI�c���5#��`e���%	f޲�:o�a�!��_��'�pM-%��By�kX�w��	C<�����b~l]S04!����H(?p�5'o5O֩�'��1�ػN�E3�c:֋[�?�F��!4�k���h�E�3��A�HF�������ؾ�]k�oK��% �q�j�_%�8O7@S����3���>���N���d�x�]�q�\}�3<��M�gy]�|�9B&9ԩ{����Yoi�ؗ�0�N*aL ���ƪ�}�Z���s�����o����h:��g �T0��:�Ф~W'�I��j��fOu��*ݡ�!ᑸp���9!,\�e$�#�ۅ�>��)�(eP��4/M
�eV�auSR ��X��uC�^��j�6���D�D����d�z겋
s`�@D�@��ހ$�K�S�Xo#c�c�p+R8�]י����\ֽ̻��rB:�yc����~� l�J?1�2�!������%���&+KE#�>��O��@b]P(�.�K�3gz>"R�~ch6�Kt�J��rlc����hiع[Gd�<Dv�#��������T�PRM�6��lcđ�w��U�p
���7��l>��ڮ�o1��׶�X�������?r�H� U�$��9uL�d�^ܾ�a/&���[�w�㬑����,w�?s�FD�g�%T��n�e�������,�( Y�IL�<�Dt��(b��Ȳ�20FN5zQ��5s^�ګ�k��-o����^��1�ݝ?��u�mH徝B�C��%��n,.���5A���� '��۹`���aS����R�ڰ������Xj��ej�O�ݸ]���]En�H�"�9؝����-�ia6a�?�r��?z�ዞ�4fu(=�ɻ4�{x���^;��Ԝ�+���{��a��`6�̇��a��Nj`{�6(����b��W��7h��o�^�Tbb#��G��	���s�$�]iE	my/�p��;LzsD	&='�;̦|�;vd2bk�#�8�d����,V,��}��gQ�A �Wox��.�Eȶ�d�r)_�������'i�譽��(�l�۬���^��r��C�ܝ=��#?��a׃�����*T�*�We�o,a&�����4���O*�>�����Li����m�Q]g��ϯ�T�o��$XwƏ�Dg�j�l�W98/g�p$�<���M�aO1 ��II�:ۅ�@�e�p��ى`�g�l�`cZ��T�v��zo������zP�!���t��J/}I���@JB�!�<<�w����}�[h��P3����g���
�}�&4n�7�Nh��pYa�.EE�2`���׸+S���Hմ��.Hm@����z����;��l�B�^������G�ўa��k����Pj,���b6[n8p��jM=��Z��
�(�p��$pExd(��D��)��>�Q�G��Z���^���)��-�@�*��lJ u�mnu<��<�N��i��}�~�.��_�@���}�R�����k/�{��ݟ�+=�"���mEO�2yD��e�w��8�tz8��_�6V0�����e�DI�/Tc��M��_������)d"B���({iSe�r(z������C�J��<B���k�Hd�Ps��O=±��Zd�����bd�Î�҃cT��Q}�v�a�l�N	hr����[�w�a)�1�����2-ao�ȳ0�9�g�����
#�������3T�r&�Jz**pGG�P"�7S�_�h4iv/����oݓ��a�F����I �#����;a�\�v�;��@�\�ɨ��F0iU�>u���>+����֟�8�h�bD�+6�����0/|��^9�O�u���ʞ��U��۲��k	r���D8��2d}�6�j�t��8{��)�$�]�It}TYhh��hF̷o��,��F5����I�!�Y�7n�3���bxzY੦�H��S�8aC��$W��gͬQ"�؋�3בh��,'��d^_=8�$���{\���R����z���.�J�9�;�z�d({�z���	4���E�=�h��.�`Π��*�l`�����	Jx,H���2蜙�������ԩ���n�%3q�9w�< �AG"۬�����a��F���Rߘvΰz��BHr Ɣ云m����v?�D�C�'�l����ИV�Wxh{s%����)�37���b�+����܅	�1�syPZ�*^t�"�JG�"�k���3�Qh�F&����[WFY!��cS2R ���e���늯��{���dx��4�D4JR �4�5��m�����B�nͱ�RAr���&F�ឱQR�~�;>��t	��`4�f;&nn�1�u��sF��aΟ��RA؎ދ�N�VE�+f�A!y�H�u,�/���}
�Z'0���ю��ޅg������9����14Z��������	_��%�D��(=�F��ug�_�*[;��� <����4Z��/i�G	]	����$���y��o�s���y~_��on�f��D΁�tf������~���ǳ�#����[H������H�b��4��!����E����_1�=��y��2�uӳE����3.�l����+l�N5O�	�sb`l���"���c����zY�K�-}��^��V��{��b]zNߜ�MsY�vc�r��fɸë�v��	����Y�#�?�ˀUgp�(??94`��< �"8m�i���t{^��i ���Y�Z�ٰb�*[o�6�e�CI�k��R��V�.���Q�[�� �
s]�,����&����Q1Q��x+_�)K�{�ǣ�=��@蠁�y[~��]l����K�N ��YE=���K����š���I�F�0y��^)�O���ajv|�(#J�u�%�Tj{�BT�gZ�*r�E�ˋ�7 �V?e��Ɇ�T�$,�9bE$٣@^�"�|ڣ��}�{�'|�����M��{�*����!-(;n����UrS���!"�aV"��>/u�o�����n�҃z�	G��&�9� ��G��ҝ?�|��XN�1_lv��/�#%o�^7ϐ������<pc�ڽ���-�~�M��O���gr���&)��I�B���^��.X1�{S�Q��33K�O�<��IDH �s��W6k�-��Ny4�I��{���TI��"�l����C�R�\�-���O�t������]i���`u��f��o�bE�n�9��DJ�Fχ;�Ł��C�Oƍ���7���૏�A��ݯ�v�v�����^�?5 <.�͸������ 
�"i��R͈�%2�ʰ�C]��Pq(O��m�&�J�լ����X�R̲U���M~j.c�pr���>:������>�M��oSw];F��g�K� :\����~'�*�\�E ��}�_�*��B��l�x���n��mr�ź��/�O�.���u�F�Og,u��	]rV��GW�T}���x��脆����B��΂�'"���� =DDl���v��ձ[��D;Q�j�.��i|�Uɰ]Q;�/q�5�7%W����R/`.H���o���I/y�E�7��> ��];<�ȭ<����K����-��@8~Kl�{�\|T����m���d��z4q�G�A�#F���.b�x�K+�^��'�~��cŇ�+D�+����s[�#�,,���.k��!*G�S�39���C�^8��,��um�Ѯ��wK;��n�<�� ':��폴����I�߿z���i�F7p6șz����G�����?��-P��WoA�2WPĐ��B�$�n���k����	����#�� �.�-灟��JpW�p�񳖜���,��XYn2��7K������ e`�L�[<�=R�:��ĐW)(����~�%�҇#(�ӈ ���#��-�<)��몮U&�Ͻ��!��P��� dD�oE}h��g��2I���W\�b��l�� �
����o��C�	��j)Z�3�<���n��U�.����w������ }��_q<`�A�����f�+�%v����^�L��'��l��{n����/&��W�Ii����}��E���`H�U�z!�� �&oy�'�-B�t{�O%PH=;�{��Z[�T��>zb���!V�cf���_��i"Aq7�,CĻ搭���a;3b��|�Y�߯�9���:-��e򻽛͒�X�t����UY/ Kӕ�Ch.I{�?'���:j�Og��g�fu
�b2�$��W��u���v2#jznA�rH������c�U5���M�X�=.�I����b�@d�Kt$#Z�mr�N�k���e%E��&j��d]y��Z=�&����o7hY��	�8�I�_�dG`�O�1��'4��o�y�5��i�O�A0^>������2f����۴N��LQR�tq�n]�)�`������l����#7��^��M�X2�'��b*po�ѫr�u�lN�"�?���D���o�o�(Z���<�H.�E|q�՟�/3�~�.dFFeN��aE�ք3E�05�4i����1Q���2��V�w ��=�DWw�,l*�2�MUA{���i۟��-�b����>�*�� J b����P�T@
�	�ёQ��d��DtrknxG�E�W[�� ^
[ňh`� N��F���Ĭ�p����^�X�������`��~kA�<\ʉ�߱��(�<[D.־r������qi�T8 ��\K|+��q���9NW&��w�ku&b��t�8�K
@��a���
����Ŕc��R���~6�B˽e J��ܠ͸w�jxF�yÈ#�	!�m�\7�5�-�P9��;�9�Z��>G���/�vGc/1>�g#�rڷqh����d,��l�0J�˳?c}à���Y�2�E����UQ�r�[�!Ve�(���؇}%AC,m1������m�[0�G2d�ͧǭ�*�!�">�Q�|�����-w�)��hy??����k�m���c�<-�AE��̆[�~�LXL$�)�ZQ~.��p��Jd������u�t�Ϧα<�n��w$��F��$�Tj]VĐ�H"aJ�3�9_��\�.�O���Ӧ�m�����;�/]�Y�4��&�i����)��<q5MJB���4����`����/;3f���瞣��!q����	�|�3��3j����'3zա�݆g��,���]�ˤŢϟ���O����L��FYLZ�om~ƆA�7�2��s�d�AM)8���/����I��$�t��*sV6�}��Kr�a��f��a���+=D*��- h׀�Lmol�K����h��-&�gs�La2WM��ٝ�����u ���c=4�{M��MTh�fw��Ȓ|!l��(���h|��,��ڣC\��Z�z�̦ a�Z��.��m��m�>|�n�p�x��f��s!)�
� 6�ک���޴��r�c��ࢮB��o�P��H�sb�w�B/��N!
�S��Y�7��t}�$��[����c{�+O=r0}�(��GS���(��>_c�&�W5�]�;�I�I[�Mz����3�*o=�b�70W��Sٰ�5�����{)�,�0B�U�����)DG*�D�.Dt�v��)0��i����̈e7���g���m}e�K$��Z�� MR���}�#/F�
�l���lz&̑���gpU�$h��<l��ф�X����f�mh�ltr���<!�G9�9OR��j�����+G.��*������%:��,D�޹*l�e-�K����Gv������Y�S�+��q[�i#�Ն��`�%Ԭ�[���iR��ʭ$Ve%f�u�qg�'�O�
n�3�Ô����f���x/��/I{ɰr%�^��`3
캴*�\�og�UpOml�+��K]U�o���)}T{.A� x���z����\=�Z�����s� ��	�Krn�┇=���_����a�҇[f]u&FD�Y��Bڞ����.�c�-��G:Pߕfy �Mt.��0%�h�;�j���n��đ�N�BC>+��Ob����T�2�����GYg��F��8<L�½�u,���b��N����]�f8M��M��#�$Nן�n|1�o�)ᔸ� x�_�S�I�Kο��f-�|$�<��["�^���/�k��z���?���?����4� 9�6���#管��By;I��e7v1)[]Gػ�N��ia�����+�_Qe�=d��(�*��31-��_b"��*62@\>�V���T�6u$̄�Ե�s�nt��Ŧk�/宎Y�6���;�6�R��/>"!X�֋�H���l�{��p�$�E�b�����T�ū6G �qV7h�4�:VhI�P���H�	|��󣄿�����sC��*<� |#��=@��=ZE��ę�Ԍ09d�Xh9}?�?�{��"{h�jL��=6�^��\��n4c��bv�3�s=o�GyLM����a��>�A����i��8Atw��pI�cͮ (�5�o
�0��XN�;X&��\���Z��k���lY�փ�TK���ǁ��9������a8��k�Gү�����g��2#��u;lb�o���ɗ�I�h���Qa�O�A��	��LdUG���a�^����͗��Dآ�&}ru���`؞7�����\��؍yv���Q��Xs�C�6
�5+�"���#\�4.��t 
����6��>1�+B[c3��>EһE�1�⛱)l��VB�)���f���V�$�/'�RL�I�)����JS�@z����H<���, �����\Y��4~�9,�nM��M��I���H�z�7ߥ�ʃd��6��D�U��w�j���Wx�(�Ko�=6W=l�����"��1��dr�	��+O�I6E�KB*(	�y���o�����K�L�j�V��孝�c�۔�X{������@�`�鏇�U_��
����+���gU����;.{�&�"ia�����=��V����~3�5�����.'���[o`��g��<�� ��9�6̶�dE�-�>�����y59a"�Tuo��mt��I0�3y��aKC�җ �a�}��"ie�x7�_�f�l��x��M��o��B)E�1�����	�R%���Ճ�P��a>�5�c�FO�/>�gC���3�!�^
h0Yq�(��3Q䤋��5?�0o�JE:_��h�Vl՜d�ݫ���a	*|s��y�;Zѓ(�v���ZB�9n�;R:Є��Ѷ-���m"H�dww[qᕬ��Z��������r5������1u�~�!�����͠9��3>ǈ6��Y%�lw�3P�<���y�C��(����FIΠ�J�/6D��	�5�;�Ęb�ru��~����$������ЇXi�u�h͏���|%DvT�1a��\}��F��e�}۾p>E#>��>�v��4(���ג��`��0�9�p��l�l�o���pL�_��vg"��K��������+w��9��]:}�G�@^��jJa�@�p���Ypan)i|�<���p��@��k"]/,4g�F�8Tժ���L�	�v
�0ПG�C= }K�Ãt�Ԕ\I�
ƕ�mJdݸ*�䩭[�\�M �ɬ�(�m;�����5}��.}�}�=�BMG���0kI�����S[���i,_OB��a\|G�c��+��U������d�JT}p�W~���v�a��I�R���M��HO,W�9����=��1>�QͪcX��!`]o#��_���l�ó�T"�t�.�������M��!̈́�������6�>'sFt"#K�Դ����;����]<�,v��Z����f��cj�˄��`�ø��~�#��6�nւ�o�a@��Y}�~�$��ן:)Z�'��E�0)�̂O��-&(%~�D�L����jl@e����̅�0m|��eM��G)J��%�v�{ҥ�:T�E�9�6�k;�$z��IP.(�Лp�غ����L�4cn�.+��h���n�����8F_O�5���l��cQrxsOقp݄��M�4;��K��Yd	^�Q�Q��3�N��n��m����������I��E4fd8�����m.8���\�Sñ�9��]�}�Yy�n#ƞ5?�tT��D#�=N��,nHݓ�!���sf=�aaj{4<n�;b�<V� ۜG�d���u�|��NOߔo���xr�-I�OD���m�y�=��pz-.�AjVng䋣i������Y�#V�5+C$O~c�@��j]�d���j���A��:��SEueN۶�� EN����mu�����!��-�K��b��R��h�g")w�?�ݚ��o��M����:s���	��}�������ڜ���W��@c��OZt�z�o�Tڥ4��g�V�9��e.w��]`���p�d�3~a:Ǧ\Z�i�Hu$�jd�<��b��q��Sc���O� dp&��ւ)�2*���C�)��>���F�`J�������7��b��I��u�}!mH���.�õX�^�z����)�>��x�Q#�L7�dO�;���ǁ�w�sV��F�]FՄ�@�d�������!#ȭ�ɺ�F��R����E��/����;!+�����A�z�R���_X߁ė �@D.[�J�&
��x�Jp��J��	.�i�m��/Lj�
;�1�������+L�g?Y�]���V�Q8ڡ1��ۥ��J�G��1L��J�l���*d� �rRZ#]���l+�tM��78���;��ў�wr�M��z�� l$��m��Pe5�C�P�\��|œ7�0�������E�	x�$����{��.��~hR7^c�B�ץy�K���+��CHQ�ܽZ�fc������l�·�]�Xs@� t�>�mfՓ��j퍞�����o{�
?���eM+.6!k�Yo�$ɝ��S�b�o�0#ƿ�?���H*(��q0ҳ� rmwe�M��>va7��&{iu����� �P��;�׏%M����ʛ��D�U�i�/w�ǚf���D������/kn�\�9�#a�->����y��@���TC�{/��N��O���X��sS�.,�q��\�_� @^vs�
[C�ך���d�4�Z:����{/����0� �IТ/z&���)75hӗ@_%D��%�9�P��.?��21��o�SG߸Ѵ^�a~ZXS�,�% ������&k�̔k}_t���������-0g@2��":_(s��ݒ�1���c�B�;m��(<a�!�t��;>.Yg����hN~%�L�R�4w<:g�������1�k�Bǘ�u��o����pQX䳶�m�/��4(EPy��{a���dO�M��#4H��1u5�[<���Ӏ4��jCE׈��I�^��)����|�G�jb_����G�N��0�8�Bk�[l�j���<ĉQ�r�������7k��K^��V��.�I�L�����B~����؋�&(~Y�� R)����p����� N\ mp�~�,���\�:l4k��IN����JG�������[ʖJ�?W�Ҭ��OxL���b���)�&��Е�`��_��JK���F(^��n4'�>y'�����3c�
 	q��{�)ABl�8�|�.[����.yk��<ԂBx4o-S[Q�چ7�J��1kQia�>�1�c��0W�[o1��&8!`�Y�ȏ��C�tF���'�>�P�D7�"-��4x���ь4��T	T�>�*�k�\���<�ݍ��΃U��ń���2>���!6~��k�j�����n��d�h��h&޺B52v�@tn@��S��kS��%�x�R�jêR
�D^YY�� �!�H�����W��x�O�Z�x��l�B~Y4]�e&�AS�L�o-X�<=��m��������Gao��I��(�p6�`����`���i��S�W3x�ꩯt�P�
Hݣ9ԥF^�:+x�=�kJ�0��rw+�2*Td�}7�ط�N1��5�?��+���P�zg>R��<��p��(�ɝ�n���F�}'i�2��	/�W7��K'P=�4J��p��wq����?@[�ӗ��hM�f�A4VЪҲK7����C�Eూ���1�hlc��cG��7��{Y%̯�$�CQ���I
n�6��j":�r�i��g�R�c�[�4�]�����[�O~�P?F��l=(?s�7 �Q�<��o�ED�#G@� ?��0o��������[S߉+Ld��.�}M�f�5F4�PD³ �8��V���{��\q5�n��+���k�"9@��t�_rSTi�r��k�+���.�����Sh{�uǃ-@ �h���N���7s򘥗�Q�#�8$7�e�� ku�ݽM�̈́c.e�m}�k����b@�0��M$���H:��->qg��</J^�m�g���V/�@ϫ'sr�-�˘�ɥ�B�ȫ�W��5H��/���V���Z��A��Wq���3�fr�_�b��;���&����	M�z#��,��1��K�'�)]���җl�_���*g>��ŞVm��!+c�83���i�ݧt�u�z����.�7�C��ɘY}�M!ċm�M$���M<!Y���ho�M����9��WPPu��.�tl��7a�0Y_<�����Ń�ˠ�V�m�؆�ϐ�n񁸙�\�y}n��>�/j���9�|Y�l��$��5�Ij��*�C��u�y�͜�μ�,�+�Fm���$��\W��ە�m>$�NQ9p��L���_�'��(Uŷ�����4�J����8s�ӥ�����3ͪ��к9c@s���
��
v���U��F�K����I�&��8X���tY8��wF�G��F���W1v �<��Y��,�%�ȶ(������e��9�#��t��ow.��#�"�D��hx���"�n����lyϴ� Z{o�9�2�v��Pk���H����%�-�?���j>���c�~l��?��Y`C֭�b�|Z�4�CYI�{l,�b� %�����\4/9�)����t�in�yc����ͼο����M���<��O�0p}>? ku����j9�s[aX���p8y�����H"���6���Ҏ��n���cG�9¯��i> h�������6g�$V�T�x���Z�F��ױ%��M���b��PnAZ~py�q}]�%d�w�(��98�]�E�%������(o[8!��E�YR�@����M�:E���p���[����m7�<��%�<w�m�w|��	&�\A�idZ߂�t"K9i1|�4H�/~����ж0���cP�闭ޝtV���#-���G��OMB%;�,��,7���.�6��Q]��N$OC8�U,�=���M����sBP�{*K��#/�=��n̔75��$Ӂc����\d�Q���g�z��N�4�9�nBB��.�r�pq�ꅳ��T�b�>�z�;R�����[G�`�(�;lb����P �A`���u]�30弖!���]�L("v&����^EX��`�d*��\\j�ROz���{������Y_2����qF���p��j;�1��!�����`᝚��H�_D����qO/�`i�YU��X�?EԵ�M��6��/�pt�����0��7C3�N�j߆��%��o����Y��n�j�H�X�4R�Iȝ�!<���r,�b�z��Im{y~�B_�;�V_���SHN�O�^�`y�+鳰�Q\��Q[��\�w��n�c�N�ޜ-z;�3�N0�'�G�6���e��B�����0'D�d>���f�u�@��z�]V��(���� �����W��g|w"���J-]�n�x{MF�L]��OU(����6]���[��7����@!}.�vػ
h]":���@!i?�\H�N��DQ���[��B�5=9���[���j�O�㿩�<�MCq��BR�z�mc�����v7��&�ӹ)*I ���
L�����JH� ��J����\x*�����KH�O6�T:E�&t���k���,:�g��BS/u �Q�CP�5�kLI��\Y��]�j,����o3՟�v�l�G�o�|�yf�����X/*(��U���	�Ŧǉe�5�M�W�,��+Wq������lc?�>,�����
��}SƱp4�#�y[��:O�����%:����i�C�hd�	1�ņ�0|���0  ?��%�iw�~�5)̑S;72�d�2��m_Wca�ܩ��U�܇z���ũ0;VQG�Y������@�#&~�"t8�K����?��o&��ﭸ�Js'�d]��23$5� n,�B�Z���c|򃠺�g�A�a��������Y\�P�4�8`��2C�|�*j��oj8�f^���N�6�{߮[gI%��3qǏ����.�����il*�Jv�F��2j�ű$�ˍ���7���x%���2C7)��?N����߷�{!Y_Ց��R^^ W�h��c���Z$֟�;o����c�O�����+���{���:�Q�`�튓}�_��#\�ɕ��
I���B�:��ȟ��G:
���L;����t��ݦ�y.��^Ã��J%o���x������haǒJ� N�ݨ:�Y2tT��h9�Q��5>&�X�m��=�58/1��F�I.�
�#$�#>l*��Kp�_w��-�A����Y��s���ͤ��S�D;>j����7�x�a~Ubj���+��d Jy���Mt��)ń:��x���%��+�Ӽ�5�o۔:lHZ�{�aX��FR�-6�OLk-z���HC�V�R��ٕR���{��l���Iy�����e-�A��߁���	���r����3{��1�?�	�5�{%�4�������|7n���d��L���(��Oz=>G��~ߪ�"h�\q�ll���v;*�J��R����^׀7\7�Lқ��u��y<x[3>���F�k�B�Hg����9Bk!#}o��d�%t0�<�e�H�Er�;_��	��q73Dp\_<c���6����i��u�P$ ��%.2j� Y�N�e�A<�\*N��哭"�
*�y��Z�~�@;l���<�G7��/G��{�˚<monwv�t5��Z��-!}K����Ɩ��Rƃ[RKSw�G�2XM�����Le
�8�y:���&�v��	ҥ�P�.jiq�WVt��(zi�4��]~Q�rkH�p;MWhD�3}TE���&��!=�n�ZBĘ׀Z���C�ܮ�z+a<9���k�}j�&���p-��wvY�CV�-�ui���*SA�O�S�8���+[u�	N������ڏ�4���~KYTh曰I9�s�6+|>�ڹ5�yz�+�L��r6�X��,I�/�E��g���ܤZ!=4uI�K��g�W����ކ���z��G
���*�{�)�� �/`��R:~c��i�G��IT:�$G rE/� �-a'�8a�T��9��l�FV	Q�ڷaN��ݣ��t*�7�`]��� �T&�����N	`��EtS�����f�H�2񅮨ļ
v�")ݏ|hg��;� �� �iz.̰��]u��8�S3�v9;���h���B��=6G=�Nvy��5W3��j��@�t�������'�4���Y�o�*7�DO�l�8X�����<��n�4K|w�:Ʉt���ܤ��*���֔�#3�X�]��.wv���=�VCї�.��0��6�^�0�fռְ����z�d����v��>���Ad�l�s��7 
wǊI\���A1�D�̅fk6�`B��3(���)m��i�v� ^�A����}`���#�\x�Oy8�Y󩂌�kQ2i�4�h��V�'#+�.Cl���G[U۴�T�hڸ��� �Ҭ���Ā�:/4
7F�%ȋS�ɭԖ3zH��1����*�7;0�5W�^9@4z��ƙ�npGM1��� AT^N�5[�{�C��!�䝅-bQ��u�a�h�M|s��z�	���z�(�ż� �Ґ x���\�^�?M&�j�'j�nPS�}��N��C�DTT��j�1�b�����3O�1�QB��h���{��d�,�q���:5�D��EE�~��:P�ɖ�M�k-����M�W��I��W�GP��v�Ɗ��)i��4��H�ax�aݦ� 2L}���Ւ���m�.�8 ���ju0p�r{�(6���2�k���[>04&��!��M�zw�"n$�v�0�ǫ/ҠP �ⲥ�f~�\�r�<j^�M,�H�]�Ӯ���}&)��=�_M��L$9bd~>��aYE
�����{�������������!_����3IM웚�Rv'ǈ�s�Dܸ�)��枵�*1��6���L��h4;c��,}{���������TAC�-����]�{	����E�S�4ќ"�s������_~��T����
�$޴��4"���ߡ6c%��5E�f�֘�G�lN�e.���Ɓ�Y��Z�T����n 
�;�D�����4��y���Ɓ}�Y�4j���M����Vފ3�#��*ܱXϣ��x9���5�S	�"���B#��x�v~��B����g*wޢ�����U��ҫ���[X��Bmk;���v	[�z�)��g�&tzH�*ǰ�����<�Ɵ�69;���pi��O������I��l�2��2���=-m��!ګ��^���I���d�-`�1n�3ؚp8�[��`�V��P�.�*������Q�5�D5�f�$�ן�<G�ӏ��3�@G�gr@�7.�#�z�z/!-��ߟ��c���ߋv���Ԛ���5�Ϳ!�Z���'����M�R��!O�[�":8������v;��܄c�ܹh��^'�,];]�j��\�(]��P<w��8y��P�fFh�COm����ۧ��������⻝>vY?:�������q������8���H�J��#6�!%��4� ��C�
��vǽ�"�ꊲ����.30�K˷��&,���
><֝!d�&����l0���	���s
�D3c���
����ܠJ�|ؽ��ѱ���C�f��
 n$���G2�&���L�s�/�c�FP٩%�P�x/;%"�J�(_���N���������L�?���U>#h*�}�xv����nEZ����:tϊ�Z�K�7ar���0X\��y�f�^q��k����
jt�.}������6V5#C��x��&�CgW��ȇ����R�T��=�%D��&�OC�M �*x���O�����9n5���a��5� j��t}T!H���=5�o2=δ��=\Q���إ ]�I�O����mb�X�4��0��D;��z����K��E���BTrS�����&3�����S����^	�՗�p�#��J�� y	3�H��LzxݐC@���